add20.sp SPICE FILE
.model nenh nmos
+ level = 2
+   vto = 0.688434   kp = 4.769e-05   gamma = 0.399818
+   phi = 0.85
+
+   cgso = 3.54e-10   cgdo = 3.54e-10
+   rsh = 70   cj = 0.000363
+   mj = 0.916   cjsw = 1.83e-10   mjsw = 0.195
+   tox = 2.15e-08   nsub = 1.79246e+16
+   nss = 3e+10   nfs = 10   tpg = 1
+   xj = 9e-07   ld = -8.3e-08   uo = 683.594
+   ucrit = 200   uexp = 0.0177713
+   vmax = 81459.2   neff = 2.18502
+
+   delta = 2.72869
.model penh pmos
+ level = 2
+   vto = -0.635779   kp = 1.91591e-05   gamma = 0.335224
+   phi = 0.85
+
+   cgso = 4.01e-10   cgdo = 4.01e-10
+   rsh = 164   cj = 0.000442
+   mj = 0.3285   cjsw = 2.34e-10   mjsw = 0.307
+   tox = 2.15e-08   nsub = 6e+17
+   nss = 3e+10   nfs = 85.3597   tpg = -1
+   xj = 1e-09   ld = -2.3e-08   uo = 41.2542
+   ucrit = 50408.2   uexp = 0.0976377
+   vmax = 42755.1   neff = 0.0107262
+
+   delta = 4.72482
m0 3 4 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.709e-11 ps=1.13e-05 pd=2.054e-05 
+ nrs=0.21 nrd=0.27 
m1 0 5 3 0 nenh l=1.1e-06 w=8e-06 
+ as=1.709e-11 ad=1.32e-11 ps=2.054e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m2 6 4 3 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m3 1 5 6 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.896e-11 ad=2.38e-11 ps=6.913e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m4 7 8 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.709e-11 ps=1.13e-05 pd=2.054e-05 
+ nrs=0.21 nrd=0.27 
m5 0 9 7 0 nenh l=1.1e-06 w=8e-06 
+ as=1.709e-11 ad=1.32e-11 ps=2.054e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m6 10 8 7 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m7 1 9 10 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.896e-11 ad=2.38e-11 ps=6.913e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m8 11 4 12 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m9 0 5 11 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.417e-11 ad=1.36e-11 ps=4.108e-05 pd=1.77e-05 
+ nrs=0.13 nrd=0.05 
m10 12 4 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.948e-11 ps=1.73e-05 pd=3.457e-05 
+ nrs=0.12 nrd=0.15 
m11 1 5 12 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.948e-11 ad=2.31e-11 ps=3.457e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m12 13 8 14 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m13 0 9 13 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.417e-11 ad=1.36e-11 ps=4.108e-05 pd=1.77e-05 
+ nrs=0.13 nrd=0.05 
m14 14 8 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.948e-11 ps=1.73e-05 pd=3.457e-05 
+ nrs=0.12 nrd=0.15 
m15 1 9 14 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.948e-11 ad=2.31e-11 ps=3.457e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m16 15 16 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.709e-11 ps=1.13e-05 pd=2.054e-05 
+ nrs=0.21 nrd=0.27 
m17 0 17 15 0 nenh l=1.1e-06 w=8e-06 
+ as=1.709e-11 ad=1.32e-11 ps=2.054e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m18 18 16 15 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m19 1 17 18 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.896e-11 ad=2.38e-11 ps=6.913e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m20 19 20 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.709e-11 ps=1.13e-05 pd=2.054e-05 
+ nrs=0.21 nrd=0.27 
m21 0 21 19 0 nenh l=1.1e-06 w=8e-06 
+ as=1.709e-11 ad=1.32e-11 ps=2.054e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m22 22 20 19 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m23 1 21 22 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.896e-11 ad=2.38e-11 ps=6.913e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m24 0 19 23 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.794e-11 ad=2.562e-11 ps=2.157e-05 pd=2.29e-05 
+ nrs=0.25 nrd=0.36 
m25 1 19 23 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.285e-11 ad=2.694e-11 ps=3.852e-05 pd=3.57e-05 
+ nrs=0.13 nrd=0.11 
m26 24 7 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.709e-11 ps=1.13e-05 pd=2.054e-05 
+ nrs=0.21 nrd=0.27 
m27 0 25 24 0 nenh l=1.1e-06 w=8e-06 
+ as=1.709e-11 ad=1.32e-11 ps=2.054e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m28 26 7 24 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m29 1 25 26 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.896e-11 ad=2.38e-11 ps=6.913e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m30 27 28 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.709e-11 ps=1.13e-05 pd=2.054e-05 
+ nrs=0.21 nrd=0.27 
m31 0 7 27 0 nenh l=1.1e-06 w=8e-06 
+ as=1.709e-11 ad=1.32e-11 ps=2.054e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m32 29 28 27 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m33 1 7 29 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.896e-11 ad=2.38e-11 ps=6.913e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m34 0 27 30 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.794e-11 ad=2.562e-11 ps=2.157e-05 pd=2.29e-05 
+ nrs=0.25 nrd=0.36 
m35 1 27 30 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.285e-11 ad=2.694e-11 ps=3.852e-05 pd=3.57e-05 
+ nrs=0.13 nrd=0.11 
m36 25 31 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.709e-11 ps=1.13e-05 pd=2.054e-05 
+ nrs=0.21 nrd=0.27 
m37 0 32 25 0 nenh l=1.1e-06 w=8e-06 
+ as=1.709e-11 ad=1.32e-11 ps=2.054e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m38 33 31 25 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m39 1 32 33 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.896e-11 ad=2.38e-11 ps=6.913e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m40 0 25 34 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.794e-11 ad=2.562e-11 ps=2.157e-05 pd=2.29e-05 
+ nrs=0.25 nrd=0.36 
m41 1 25 34 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.285e-11 ad=2.694e-11 ps=3.852e-05 pd=3.57e-05 
+ nrs=0.13 nrd=0.11 
m42 35 36 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.709e-11 ps=1.13e-05 pd=2.054e-05 
+ nrs=0.21 nrd=0.27 
m43 0 37 35 0 nenh l=1.1e-06 w=8e-06 
+ as=1.709e-11 ad=1.32e-11 ps=2.054e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m44 38 36 35 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m45 1 37 38 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.896e-11 ad=2.38e-11 ps=6.913e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m46 39 40 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.709e-11 ps=1.13e-05 pd=2.054e-05 
+ nrs=0.21 nrd=0.27 
m47 0 41 39 0 nenh l=1.1e-06 w=8e-06 
+ as=1.709e-11 ad=1.32e-11 ps=2.054e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m48 42 40 39 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m49 1 41 42 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.896e-11 ad=2.38e-11 ps=6.913e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m50 43 30 44 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m51 0 14 43 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.417e-11 ad=1.36e-11 ps=4.108e-05 pd=1.77e-05 
+ nrs=0.13 nrd=0.05 
m52 44 30 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.948e-11 ps=1.73e-05 pd=3.457e-05 
+ nrs=0.12 nrd=0.15 
m53 1 14 44 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.948e-11 ad=2.31e-11 ps=3.457e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m54 45 16 46 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m55 0 17 45 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.417e-11 ad=1.36e-11 ps=4.108e-05 pd=1.77e-05 
+ nrs=0.13 nrd=0.05 
m56 46 16 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.948e-11 ps=1.73e-05 pd=3.457e-05 
+ nrs=0.12 nrd=0.15 
m57 1 17 46 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.948e-11 ad=2.31e-11 ps=3.457e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m58 47 24 48 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m59 0 23 47 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.417e-11 ad=1.36e-11 ps=4.108e-05 pd=1.77e-05 
+ nrs=0.13 nrd=0.05 
m60 48 24 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.948e-11 ps=1.73e-05 pd=3.457e-05 
+ nrs=0.12 nrd=0.15 
m61 1 23 48 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.948e-11 ad=2.31e-11 ps=3.457e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m62 49 20 50 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m63 0 21 49 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.417e-11 ad=1.36e-11 ps=4.108e-05 pd=1.77e-05 
+ nrs=0.13 nrd=0.05 
m64 50 20 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.948e-11 ps=1.73e-05 pd=3.457e-05 
+ nrs=0.12 nrd=0.15 
m65 1 21 50 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.948e-11 ad=2.31e-11 ps=3.457e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m66 51 31 28 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m67 0 32 51 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.417e-11 ad=1.36e-11 ps=4.108e-05 pd=1.77e-05 
+ nrs=0.13 nrd=0.05 
m68 28 31 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.948e-11 ps=1.73e-05 pd=3.457e-05 
+ nrs=0.12 nrd=0.15 
m69 1 32 28 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.948e-11 ad=2.31e-11 ps=3.457e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m70 52 36 53 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m71 0 37 52 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.417e-11 ad=1.36e-11 ps=4.108e-05 pd=1.77e-05 
+ nrs=0.13 nrd=0.05 
m72 53 36 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.948e-11 ps=1.73e-05 pd=3.457e-05 
+ nrs=0.12 nrd=0.15 
m73 1 37 53 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.948e-11 ad=2.31e-11 ps=3.457e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m74 54 40 55 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m75 0 41 54 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.417e-11 ad=1.36e-11 ps=4.108e-05 pd=1.77e-05 
+ nrs=0.13 nrd=0.05 
m76 55 40 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.948e-11 ps=1.73e-05 pd=3.457e-05 
+ nrs=0.12 nrd=0.15 
m77 1 41 55 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.948e-11 ad=2.31e-11 ps=3.457e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m78 56 46 57 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m79 0 58 56 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.417e-11 ad=2.507e-11 ps=4.108e-05 pd=2.557e-05 
+ nrs=0.13 nrd=0.1 
m80 56 15 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.417e-11 ps=2.557e-05 pd=4.108e-05 
+ nrs=0.1 nrd=0.13 
m81 57 46 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.896e-11 ps=3.13e-05 pd=6.913e-05 
+ nrs=0.06 nrd=0.08 
m82 59 58 57 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m83 1 15 59 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.896e-11 ad=4.62e-11 ps=6.913e-05 pd=3.13e-05 
+ nrs=0.08 nrd=0.06 
m84 0 15 60 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.794e-11 ad=2.562e-11 ps=2.157e-05 pd=2.29e-05 
+ nrs=0.25 nrd=0.36 
m85 1 15 60 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.285e-11 ad=2.694e-11 ps=3.852e-05 pd=3.57e-05 
+ nrs=0.13 nrd=0.11 
m86 58 61 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.709e-11 ps=1.13e-05 pd=2.054e-05 
+ nrs=0.21 nrd=0.27 
m87 0 62 58 0 nenh l=1.1e-06 w=8e-06 
+ as=1.709e-11 ad=1.32e-11 ps=2.054e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m88 63 61 58 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m89 1 62 63 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.896e-11 ad=2.38e-11 ps=6.913e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m90 0 58 64 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.794e-11 ad=2.562e-11 ps=2.157e-05 pd=2.29e-05 
+ nrs=0.25 nrd=0.36 
m91 1 58 64 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.285e-11 ad=2.694e-11 ps=3.852e-05 pd=3.57e-05 
+ nrs=0.13 nrd=0.11 
m92 65 53 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.709e-11 ps=1.13e-05 pd=2.054e-05 
+ nrs=0.21 nrd=0.27 
m93 0 39 65 0 nenh l=1.1e-06 w=8e-06 
+ as=1.709e-11 ad=1.32e-11 ps=2.054e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m94 66 53 65 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m95 1 39 66 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.896e-11 ad=2.38e-11 ps=6.913e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m96 0 55 67 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.794e-11 ad=2.562e-11 ps=2.157e-05 pd=2.29e-05 
+ nrs=0.25 nrd=0.36 
m97 1 55 67 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.285e-11 ad=2.694e-11 ps=3.852e-05 pd=3.57e-05 
+ nrs=0.13 nrd=0.11 
m98 68 67 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.709e-11 ps=1.13e-05 pd=2.054e-05 
+ nrs=0.21 nrd=0.27 
m99 0 39 68 0 nenh l=1.1e-06 w=8e-06 
+ as=1.709e-11 ad=1.32e-11 ps=2.054e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m100 69 67 68 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m101 1 39 69 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.896e-11 ad=2.38e-11 ps=6.913e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m102 70 71 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.709e-11 ps=1.13e-05 pd=2.054e-05 
+ nrs=0.21 nrd=0.27 
m103 0 72 70 0 nenh l=1.1e-06 w=8e-06 
+ as=1.709e-11 ad=1.32e-11 ps=2.054e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m104 73 71 70 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m105 1 72 73 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.896e-11 ad=2.38e-11 ps=6.913e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m106 74 46 75 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m107 0 60 74 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.417e-11 ad=1.36e-11 ps=4.108e-05 pd=1.77e-05 
+ nrs=0.13 nrd=0.05 
m108 75 46 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.948e-11 ps=1.73e-05 pd=3.457e-05 
+ nrs=0.12 nrd=0.15 
m109 1 60 75 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.948e-11 ad=2.31e-11 ps=3.457e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m110 0 39 76 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.417e-11 ad=3.008e-11 ps=4.108e-05 pd=3.81e-05 
+ nrs=0.13 nrd=0.12 
m111 77 78 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=3.417e-11 ps=1.77e-05 pd=4.108e-05 
+ nrs=0.05 nrd=0.13 
m112 76 55 77 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.008e-11 ad=1.36e-11 ps=3.81e-05 pd=1.77e-05 
+ nrs=0.12 nrd=0.05 
m113 79 39 76 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=3.5e-11 ps=4.183e-05 pd=6.21e-05 
+ nrs=0.06 nrd=0.04 
m114 1 78 79 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.896e-11 ad=4.62e-11 ps=6.913e-05 pd=4.183e-05 
+ nrs=0.08 nrd=0.06 
m115 79 55 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.896e-11 ps=4.183e-05 pd=6.913e-05 
+ nrs=0.06 nrd=0.08 
m116 80 81 61 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m117 0 55 80 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.417e-11 ad=1.36e-11 ps=4.108e-05 pd=1.77e-05 
+ nrs=0.13 nrd=0.05 
m118 61 81 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.948e-11 ps=1.73e-05 pd=3.457e-05 
+ nrs=0.12 nrd=0.15 
m119 1 55 61 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.948e-11 ad=2.31e-11 ps=3.457e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m120 82 71 83 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m121 0 72 82 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.417e-11 ad=1.36e-11 ps=4.108e-05 pd=1.77e-05 
+ nrs=0.13 nrd=0.05 
m122 83 71 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.948e-11 ps=1.73e-05 pd=3.457e-05 
+ nrs=0.12 nrd=0.15 
m123 1 72 83 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.948e-11 ad=2.31e-11 ps=3.457e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m124 84 85 78 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m125 0 86 84 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.417e-11 ad=2.507e-11 ps=4.108e-05 pd=2.557e-05 
+ nrs=0.13 nrd=0.1 
m126 84 87 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.417e-11 ps=2.557e-05 pd=4.108e-05 
+ nrs=0.1 nrd=0.13 
m127 78 85 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.896e-11 ps=3.13e-05 pd=6.913e-05 
+ nrs=0.06 nrd=0.08 
m128 88 86 78 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m129 1 87 88 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.896e-11 ad=4.62e-11 ps=6.913e-05 pd=3.13e-05 
+ nrs=0.08 nrd=0.06 
m130 0 90 89 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.417e-11 ad=3.008e-11 ps=4.108e-05 pd=3.81e-05 
+ nrs=0.13 nrd=0.12 
m131 91 78 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=3.417e-11 ps=1.77e-05 pd=4.108e-05 
+ nrs=0.05 nrd=0.13 
m132 89 68 91 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.008e-11 ad=1.36e-11 ps=3.81e-05 pd=1.77e-05 
+ nrs=0.12 nrd=0.05 
m133 92 90 89 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=3.5e-11 ps=4.183e-05 pd=6.21e-05 
+ nrs=0.06 nrd=0.04 
m134 1 78 92 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.896e-11 ad=4.62e-11 ps=6.913e-05 pd=4.183e-05 
+ nrs=0.08 nrd=0.06 
m135 92 68 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.896e-11 ps=4.183e-05 pd=6.913e-05 
+ nrs=0.06 nrd=0.08 
m136 0 68 90 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.417e-11 ad=3.008e-11 ps=4.108e-05 pd=3.81e-05 
+ nrs=0.13 nrd=0.12 
m137 93 94 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=3.417e-11 ps=1.77e-05 pd=4.108e-05 
+ nrs=0.05 nrd=0.13 
m138 90 53 93 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.008e-11 ad=1.36e-11 ps=3.81e-05 pd=1.77e-05 
+ nrs=0.12 nrd=0.05 
m139 95 68 90 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=3.5e-11 ps=4.183e-05 pd=6.21e-05 
+ nrs=0.06 nrd=0.04 
m140 1 94 95 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.896e-11 ad=4.62e-11 ps=6.913e-05 pd=4.183e-05 
+ nrs=0.08 nrd=0.06 
m141 95 53 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.896e-11 ps=4.183e-05 pd=6.913e-05 
+ nrs=0.06 nrd=0.08 
m142 0 89 96 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.794e-11 ad=2.562e-11 ps=2.157e-05 pd=2.29e-05 
+ nrs=0.25 nrd=0.36 
m143 1 89 96 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.285e-11 ad=2.694e-11 ps=3.852e-05 pd=3.57e-05 
+ nrs=0.13 nrd=0.11 
m144 0 53 87 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.794e-11 ad=2.562e-11 ps=2.157e-05 pd=2.29e-05 
+ nrs=0.25 nrd=0.36 
m145 1 53 87 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.285e-11 ad=2.694e-11 ps=3.852e-05 pd=3.57e-05 
+ nrs=0.13 nrd=0.11 
m146 97 98 94 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m147 0 85 97 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.417e-11 ad=1.36e-11 ps=4.108e-05 pd=1.77e-05 
+ nrs=0.13 nrd=0.05 
m148 94 98 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.948e-11 ps=1.73e-05 pd=3.457e-05 
+ nrs=0.12 nrd=0.15 
m149 1 85 94 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.948e-11 ad=2.31e-11 ps=3.457e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m150 99 53 100 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m151 0 85 99 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.417e-11 ad=1.36e-11 ps=4.108e-05 pd=1.77e-05 
+ nrs=0.13 nrd=0.05 
m152 100 53 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.948e-11 ps=1.73e-05 pd=3.457e-05 
+ nrs=0.12 nrd=0.15 
m153 1 85 100 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.948e-11 ad=2.31e-11 ps=3.457e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m154 101 44 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.788e-11 ps=1.13e-05 pd=1.959e-05 
+ nrs=0.21 nrd=0.28 
m155 0 102 101 0 nenh l=1.1e-06 w=8e-06 
+ as=1.788e-11 ad=1.32e-11 ps=1.959e-05 pd=1.13e-05 
+ nrs=0.28 nrd=0.21 
m156 103 44 101 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m157 1 102 103 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.054e-11 ad=2.38e-11 ps=6.96e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m158 0 104 102 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.877e-11 ad=2.562e-11 ps=2.057e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m159 1 104 102 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.373e-11 ad=2.694e-11 ps=3.878e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m160 0 3 105 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.877e-11 ad=2.562e-11 ps=2.057e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m161 1 3 105 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.373e-11 ad=2.694e-11 ps=3.878e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m162 0 14 106 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.877e-11 ad=2.562e-11 ps=2.057e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m163 1 14 106 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.373e-11 ad=2.694e-11 ps=3.878e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m164 107 106 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.788e-11 ps=1.13e-05 pd=1.959e-05 
+ nrs=0.21 nrd=0.28 
m165 0 7 107 0 nenh l=1.1e-06 w=8e-06 
+ as=1.788e-11 ad=1.32e-11 ps=1.959e-05 pd=1.13e-05 
+ nrs=0.28 nrd=0.21 
m166 108 106 107 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m167 1 7 108 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.054e-11 ad=2.38e-11 ps=6.96e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m168 109 110 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.788e-11 ps=1.13e-05 pd=1.959e-05 
+ nrs=0.21 nrd=0.28 
m169 0 111 109 0 nenh l=1.1e-06 w=8e-06 
+ as=1.788e-11 ad=1.32e-11 ps=1.959e-05 pd=1.13e-05 
+ nrs=0.28 nrd=0.21 
m170 112 110 109 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m171 1 111 112 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.054e-11 ad=2.38e-11 ps=6.96e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m172 0 114 113 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.877e-11 ad=2.562e-11 ps=2.057e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m173 1 114 113 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.373e-11 ad=2.694e-11 ps=3.878e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m174 115 116 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.788e-11 ps=1.13e-05 pd=1.959e-05 
+ nrs=0.21 nrd=0.28 
m175 0 19 115 0 nenh l=1.1e-06 w=8e-06 
+ as=1.788e-11 ad=1.32e-11 ps=1.959e-05 pd=1.13e-05 
+ nrs=0.28 nrd=0.21 
m176 117 116 115 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m177 1 19 117 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.054e-11 ad=2.38e-11 ps=6.96e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m178 0 50 116 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.877e-11 ad=2.562e-11 ps=2.057e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m179 1 50 116 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.373e-11 ad=2.694e-11 ps=3.878e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m180 118 24 104 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m181 0 116 118 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.575e-11 ad=1.36e-11 ps=3.918e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m182 104 24 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=3.027e-11 ps=1.73e-05 pd=3.48e-05 
+ nrs=0.12 nrd=0.15 
m183 1 116 104 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.027e-11 ad=2.31e-11 ps=3.48e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m184 0 7 119 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.575e-11 ad=3.008e-11 ps=3.918e-05 pd=3.81e-05 
+ nrs=0.14 nrd=0.12 
m185 120 121 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=3.575e-11 ps=1.77e-05 pd=3.918e-05 
+ nrs=0.05 nrd=0.14 
m186 119 14 120 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.008e-11 ad=1.36e-11 ps=3.81e-05 pd=1.77e-05 
+ nrs=0.12 nrd=0.05 
m187 122 7 119 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=3.5e-11 ps=4.183e-05 pd=6.21e-05 
+ nrs=0.06 nrd=0.04 
m188 1 121 122 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.054e-11 ad=4.62e-11 ps=6.96e-05 pd=4.183e-05 
+ nrs=0.08 nrd=0.06 
m189 122 14 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=6.054e-11 ps=4.183e-05 pd=6.96e-05 
+ nrs=0.06 nrd=0.08 
m190 123 110 114 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m191 0 111 123 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.575e-11 ad=1.36e-11 ps=3.918e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m192 114 110 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=3.027e-11 ps=1.73e-05 pd=3.48e-05 
+ nrs=0.12 nrd=0.15 
m193 1 111 114 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.027e-11 ad=2.31e-11 ps=3.48e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m194 0 125 124 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.575e-11 ad=3.008e-11 ps=3.918e-05 pd=3.81e-05 
+ nrs=0.14 nrd=0.12 
m195 126 121 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=3.575e-11 ps=1.77e-05 pd=3.918e-05 
+ nrs=0.05 nrd=0.14 
m196 124 107 126 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.008e-11 ad=1.36e-11 ps=3.81e-05 pd=1.77e-05 
+ nrs=0.12 nrd=0.05 
m197 127 125 124 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=3.5e-11 ps=4.183e-05 pd=6.21e-05 
+ nrs=0.06 nrd=0.04 
m198 1 121 127 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.054e-11 ad=4.62e-11 ps=6.96e-05 pd=4.183e-05 
+ nrs=0.08 nrd=0.06 
m199 127 107 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=6.054e-11 ps=4.183e-05 pd=6.96e-05 
+ nrs=0.06 nrd=0.08 
m200 0 107 125 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.575e-11 ad=3.008e-11 ps=3.918e-05 pd=3.81e-05 
+ nrs=0.14 nrd=0.12 
m201 128 129 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=3.575e-11 ps=1.77e-05 pd=3.918e-05 
+ nrs=0.05 nrd=0.14 
m202 125 28 128 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.008e-11 ad=1.36e-11 ps=3.81e-05 pd=1.77e-05 
+ nrs=0.12 nrd=0.05 
m203 130 107 125 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=3.5e-11 ps=4.183e-05 pd=6.21e-05 
+ nrs=0.06 nrd=0.04 
m204 1 129 130 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.054e-11 ad=4.62e-11 ps=6.96e-05 pd=4.183e-05 
+ nrs=0.08 nrd=0.06 
m205 130 28 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=6.054e-11 ps=4.183e-05 pd=6.96e-05 
+ nrs=0.06 nrd=0.08 
m206 131 132 129 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m207 0 34 131 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.575e-11 ad=1.36e-11 ps=3.918e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m208 129 132 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=3.027e-11 ps=1.73e-05 pd=3.48e-05 
+ nrs=0.12 nrd=0.15 
m209 1 34 129 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.027e-11 ad=2.31e-11 ps=3.48e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m210 0 28 133 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.877e-11 ad=2.562e-11 ps=2.057e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m211 1 28 133 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.373e-11 ad=2.694e-11 ps=3.878e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m212 134 28 135 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m213 0 34 134 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.575e-11 ad=1.36e-11 ps=3.918e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m214 135 28 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=3.027e-11 ps=1.73e-05 pd=3.48e-05 
+ nrs=0.12 nrd=0.15 
m215 1 34 135 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.027e-11 ad=2.31e-11 ps=3.48e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m216 136 34 121 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m217 0 137 136 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.575e-11 ad=2.507e-11 ps=3.918e-05 pd=2.557e-05 
+ nrs=0.14 nrd=0.1 
m218 136 133 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.575e-11 ps=2.557e-05 pd=3.918e-05 
+ nrs=0.1 nrd=0.14 
m219 121 34 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=6.054e-11 ps=3.13e-05 pd=6.96e-05 
+ nrs=0.06 nrd=0.08 
m220 138 137 121 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m221 1 133 138 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.054e-11 ad=4.62e-11 ps=6.96e-05 pd=3.13e-05 
+ nrs=0.08 nrd=0.06 
m222 0 109 139 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.877e-11 ad=2.562e-11 ps=2.057e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m223 1 109 139 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.373e-11 ad=2.694e-11 ps=3.878e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m224 140 39 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.788e-11 ps=1.13e-05 pd=1.959e-05 
+ nrs=0.21 nrd=0.28 
m225 0 35 140 0 nenh l=1.1e-06 w=8e-06 
+ as=1.788e-11 ad=1.32e-11 ps=1.959e-05 pd=1.13e-05 
+ nrs=0.28 nrd=0.21 
m226 141 39 140 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m227 1 35 141 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.054e-11 ad=2.38e-11 ps=6.96e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m228 0 142 62 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.877e-11 ad=2.562e-11 ps=2.057e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m229 1 142 62 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.373e-11 ad=2.694e-11 ps=3.878e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m230 0 35 85 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.877e-11 ad=2.562e-11 ps=2.057e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m231 1 35 85 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.373e-11 ad=2.694e-11 ps=3.878e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m232 143 144 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.788e-11 ps=1.13e-05 pd=1.959e-05 
+ nrs=0.21 nrd=0.28 
m233 0 145 143 0 nenh l=1.1e-06 w=8e-06 
+ as=1.788e-11 ad=1.32e-11 ps=1.959e-05 pd=1.13e-05 
+ nrs=0.28 nrd=0.21 
m234 146 144 143 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m235 1 145 146 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.054e-11 ad=2.38e-11 ps=6.96e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m236 147 140 142 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m237 0 113 147 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.575e-11 ad=1.36e-11 ps=3.918e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m238 142 140 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=3.027e-11 ps=1.73e-05 pd=3.48e-05 
+ nrs=0.12 nrd=0.15 
m239 1 113 142 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.027e-11 ad=2.31e-11 ps=3.48e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m240 148 144 149 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m241 0 145 148 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.575e-11 ad=1.36e-11 ps=3.918e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m242 149 144 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=3.027e-11 ps=1.73e-05 pd=3.48e-05 
+ nrs=0.12 nrd=0.15 
m243 1 145 149 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.027e-11 ad=2.31e-11 ps=3.48e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m244 150 152 151 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m245 0 76 150 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.575e-11 ad=2.507e-11 ps=3.918e-05 pd=2.557e-05 
+ nrs=0.14 nrd=0.1 
m246 150 75 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.575e-11 ps=2.557e-05 pd=3.918e-05 
+ nrs=0.1 nrd=0.14 
m247 151 152 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=6.054e-11 ps=3.13e-05 pd=6.96e-05 
+ nrs=0.06 nrd=0.08 
m248 153 76 151 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m249 1 75 153 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.054e-11 ad=4.62e-11 ps=6.96e-05 pd=3.13e-05 
+ nrs=0.08 nrd=0.06 
m250 154 75 152 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m251 0 155 154 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.575e-11 ad=2.507e-11 ps=3.918e-05 pd=2.557e-05 
+ nrs=0.14 nrd=0.1 
m252 154 64 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.575e-11 ps=2.557e-05 pd=3.918e-05 
+ nrs=0.1 nrd=0.14 
m253 152 75 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=6.054e-11 ps=3.13e-05 pd=6.96e-05 
+ nrs=0.06 nrd=0.08 
m254 156 155 152 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m255 1 64 156 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.054e-11 ad=4.62e-11 ps=6.96e-05 pd=3.13e-05 
+ nrs=0.08 nrd=0.06 
m256 157 158 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.788e-11 ps=1.13e-05 pd=1.959e-05 
+ nrs=0.21 nrd=0.28 
m257 0 159 157 0 nenh l=1.1e-06 w=8e-06 
+ as=1.788e-11 ad=1.32e-11 ps=1.959e-05 pd=1.13e-05 
+ nrs=0.28 nrd=0.21 
m258 160 158 157 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m259 1 159 160 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.054e-11 ad=2.38e-11 ps=6.96e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m260 0 157 161 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.877e-11 ad=2.562e-11 ps=2.057e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m261 1 157 161 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.373e-11 ad=2.694e-11 ps=3.878e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m262 0 65 81 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.877e-11 ad=2.562e-11 ps=2.057e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m263 1 65 81 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.373e-11 ad=2.694e-11 ps=3.878e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m264 162 163 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.788e-11 ps=1.13e-05 pd=1.959e-05 
+ nrs=0.21 nrd=0.28 
m265 0 164 162 0 nenh l=1.1e-06 w=8e-06 
+ as=1.788e-11 ad=1.32e-11 ps=1.959e-05 pd=1.13e-05 
+ nrs=0.28 nrd=0.21 
m266 165 163 162 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m267 1 164 165 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.054e-11 ad=2.38e-11 ps=6.96e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m268 166 109 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.788e-11 ps=1.13e-05 pd=1.959e-05 
+ nrs=0.21 nrd=0.28 
m269 0 167 166 0 nenh l=1.1e-06 w=8e-06 
+ as=1.788e-11 ad=1.32e-11 ps=1.959e-05 pd=1.13e-05 
+ nrs=0.28 nrd=0.21 
m270 168 109 166 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m271 1 167 168 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.054e-11 ad=2.38e-11 ps=6.96e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m272 0 170 169 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.877e-11 ad=2.562e-11 ps=2.057e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m273 1 170 169 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.373e-11 ad=2.694e-11 ps=3.878e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m274 0 166 171 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.877e-11 ad=2.562e-11 ps=2.057e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m275 1 166 171 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.373e-11 ad=2.694e-11 ps=3.878e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m276 172 158 173 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m277 0 159 172 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.575e-11 ad=1.36e-11 ps=3.918e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m278 173 158 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=3.027e-11 ps=1.73e-05 pd=3.48e-05 
+ nrs=0.12 nrd=0.15 
m279 1 159 173 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.027e-11 ad=2.31e-11 ps=3.48e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m280 174 163 175 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m281 0 164 174 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.575e-11 ad=1.36e-11 ps=3.918e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m282 175 163 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=3.027e-11 ps=1.73e-05 pd=3.48e-05 
+ nrs=0.12 nrd=0.15 
m283 1 164 175 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.027e-11 ad=2.31e-11 ps=3.48e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m284 176 114 170 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m285 0 167 176 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.575e-11 ad=1.36e-11 ps=3.918e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m286 170 114 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=3.027e-11 ps=1.73e-05 pd=3.48e-05 
+ nrs=0.12 nrd=0.15 
m287 1 167 170 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.027e-11 ad=2.31e-11 ps=3.48e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m288 177 171 98 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m289 0 114 177 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.575e-11 ad=1.36e-11 ps=3.918e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m290 98 171 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=3.027e-11 ps=1.73e-05 pd=3.48e-05 
+ nrs=0.12 nrd=0.15 
m291 1 114 98 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.027e-11 ad=2.31e-11 ps=3.48e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m292 178 173 179 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m293 0 161 178 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.575e-11 ad=1.36e-11 ps=3.918e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m294 179 173 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=3.027e-11 ps=1.73e-05 pd=3.48e-05 
+ nrs=0.12 nrd=0.15 
m295 1 161 179 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.027e-11 ad=2.31e-11 ps=3.48e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m296 180 182 181 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m297 0 161 180 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.575e-11 ad=1.36e-11 ps=3.918e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m298 181 182 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=3.027e-11 ps=1.73e-05 pd=3.48e-05 
+ nrs=0.12 nrd=0.15 
m299 1 161 181 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.027e-11 ad=2.31e-11 ps=3.48e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m300 183 161 184 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m301 0 185 183 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.575e-11 ad=2.507e-11 ps=3.918e-05 pd=2.557e-05 
+ nrs=0.14 nrd=0.1 
m302 183 186 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.575e-11 ps=2.557e-05 pd=3.918e-05 
+ nrs=0.1 nrd=0.14 
m303 184 161 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=6.054e-11 ps=3.13e-05 pd=6.96e-05 
+ nrs=0.06 nrd=0.08 
m304 187 185 184 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m305 1 186 187 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.054e-11 ad=4.62e-11 ps=6.96e-05 pd=3.13e-05 
+ nrs=0.08 nrd=0.06 
m306 0 101 188 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.806e-11 ad=2.562e-11 ps=2.064e-05 pd=2.29e-05 
+ nrs=0.26 nrd=0.36 
m307 1 101 188 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.211e-11 ad=2.694e-11 ps=3.927e-05 pd=3.57e-05 
+ nrs=0.13 nrd=0.11 
m308 189 48 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.72e-11 ps=1.13e-05 pd=1.966e-05 
+ nrs=0.21 nrd=0.27 
m309 0 3 189 0 nenh l=1.1e-06 w=8e-06 
+ as=1.72e-11 ad=1.32e-11 ps=1.966e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m310 190 48 189 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m311 1 3 190 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.764e-11 ad=2.38e-11 ps=7.049e-05 pd=2.97e-05 
+ nrs=0.07 nrd=0.03 
m312 191 193 192 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m313 0 189 191 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.44e-11 ad=1.36e-11 ps=3.932e-05 pd=1.77e-05 
+ nrs=0.13 nrd=0.05 
m314 192 193 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.882e-11 ps=1.73e-05 pd=3.524e-05 
+ nrs=0.12 nrd=0.15 
m315 1 189 192 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.882e-11 ad=2.31e-11 ps=3.524e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m316 194 12 195 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m317 0 105 194 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.44e-11 ad=1.36e-11 ps=3.932e-05 pd=1.77e-05 
+ nrs=0.13 nrd=0.05 
m318 195 12 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.882e-11 ps=1.73e-05 pd=3.524e-05 
+ nrs=0.12 nrd=0.15 
m319 1 105 195 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.882e-11 ad=2.31e-11 ps=3.524e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m320 196 195 197 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m321 0 198 196 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.44e-11 ad=2.507e-11 ps=3.932e-05 pd=2.557e-05 
+ nrs=0.13 nrd=0.1 
m322 196 188 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.44e-11 ps=2.557e-05 pd=3.932e-05 
+ nrs=0.1 nrd=0.13 
m323 197 195 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.764e-11 ps=3.13e-05 pd=7.049e-05 
+ nrs=0.06 nrd=0.07 
m324 199 198 197 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m325 1 188 199 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.764e-11 ad=4.62e-11 ps=7.049e-05 pd=3.13e-05 
+ nrs=0.07 nrd=0.06 
m326 200 197 201 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m327 0 119 200 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.44e-11 ad=2.507e-11 ps=3.932e-05 pd=2.557e-05 
+ nrs=0.13 nrd=0.1 
m328 200 195 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.44e-11 ps=2.557e-05 pd=3.932e-05 
+ nrs=0.1 nrd=0.13 
m329 201 197 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.764e-11 ps=3.13e-05 pd=7.049e-05 
+ nrs=0.06 nrd=0.07 
m330 202 119 201 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m331 1 195 202 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.764e-11 ad=4.62e-11 ps=7.049e-05 pd=3.13e-05 
+ nrs=0.07 nrd=0.06 
m332 198 48 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.72e-11 ps=1.13e-05 pd=1.966e-05 
+ nrs=0.21 nrd=0.27 
m333 0 203 198 0 nenh l=1.1e-06 w=8e-06 
+ as=1.72e-11 ad=1.32e-11 ps=1.966e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m334 204 48 198 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m335 1 203 204 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.764e-11 ad=2.38e-11 ps=7.049e-05 pd=2.97e-05 
+ nrs=0.07 nrd=0.03 
m336 0 193 203 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.806e-11 ad=2.562e-11 ps=2.064e-05 pd=2.29e-05 
+ nrs=0.26 nrd=0.36 
m337 1 193 203 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.211e-11 ad=2.694e-11 ps=3.927e-05 pd=3.57e-05 
+ nrs=0.13 nrd=0.11 
m338 205 207 206 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m339 0 115 205 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.44e-11 ad=2.507e-11 ps=3.932e-05 pd=2.557e-05 
+ nrs=0.13 nrd=0.1 
m340 205 203 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.44e-11 ps=2.557e-05 pd=3.932e-05 
+ nrs=0.1 nrd=0.13 
m341 206 207 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.764e-11 ps=3.13e-05 pd=7.049e-05 
+ nrs=0.06 nrd=0.07 
m342 208 115 206 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m343 1 203 208 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.764e-11 ad=4.62e-11 ps=7.049e-05 pd=3.13e-05 
+ nrs=0.07 nrd=0.06 
m344 209 115 207 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m345 0 203 209 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.44e-11 ad=1.36e-11 ps=3.932e-05 pd=1.77e-05 
+ nrs=0.13 nrd=0.05 
m346 207 115 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.882e-11 ps=1.73e-05 pd=3.524e-05 
+ nrs=0.12 nrd=0.15 
m347 1 203 207 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.882e-11 ad=2.31e-11 ps=3.524e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m348 210 19 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.72e-11 ps=1.13e-05 pd=1.966e-05 
+ nrs=0.21 nrd=0.27 
m349 0 203 210 0 nenh l=1.1e-06 w=8e-06 
+ as=1.72e-11 ad=1.32e-11 ps=1.966e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m350 211 19 210 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m351 1 203 211 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.764e-11 ad=2.38e-11 ps=7.049e-05 pd=2.97e-05 
+ nrs=0.07 nrd=0.03 
m352 0 210 212 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.806e-11 ad=2.562e-11 ps=2.064e-05 pd=2.29e-05 
+ nrs=0.26 nrd=0.36 
m353 1 210 212 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.211e-11 ad=2.694e-11 ps=3.927e-05 pd=3.57e-05 
+ nrs=0.13 nrd=0.11 
m354 213 50 214 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m355 0 203 213 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.44e-11 ad=1.36e-11 ps=3.932e-05 pd=1.77e-05 
+ nrs=0.13 nrd=0.05 
m356 214 50 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.882e-11 ps=1.73e-05 pd=3.524e-05 
+ nrs=0.12 nrd=0.15 
m357 1 203 214 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.882e-11 ad=2.31e-11 ps=3.524e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m358 215 212 132 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m359 0 50 215 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.44e-11 ad=1.36e-11 ps=3.932e-05 pd=1.77e-05 
+ nrs=0.13 nrd=0.05 
m360 132 212 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.882e-11 ps=1.73e-05 pd=3.524e-05 
+ nrs=0.12 nrd=0.15 
m361 1 50 132 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.882e-11 ad=2.31e-11 ps=3.524e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m362 216 132 217 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m363 0 135 216 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.44e-11 ad=1.36e-11 ps=3.932e-05 pd=1.77e-05 
+ nrs=0.13 nrd=0.05 
m364 217 132 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.882e-11 ps=1.73e-05 pd=3.524e-05 
+ nrs=0.12 nrd=0.15 
m365 1 135 217 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.882e-11 ad=2.31e-11 ps=3.524e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m366 218 217 219 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m367 0 137 218 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.44e-11 ad=2.507e-11 ps=3.932e-05 pd=2.557e-05 
+ nrs=0.13 nrd=0.1 
m368 218 135 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.44e-11 ps=2.557e-05 pd=3.932e-05 
+ nrs=0.1 nrd=0.13 
m369 219 217 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.764e-11 ps=3.13e-05 pd=7.049e-05 
+ nrs=0.06 nrd=0.07 
m370 220 137 219 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m371 1 135 220 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.764e-11 ad=4.62e-11 ps=7.049e-05 pd=3.13e-05 
+ nrs=0.07 nrd=0.06 
m372 137 221 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.72e-11 ps=1.13e-05 pd=1.966e-05 
+ nrs=0.21 nrd=0.27 
m373 0 19 137 0 nenh l=1.1e-06 w=8e-06 
+ as=1.72e-11 ad=1.32e-11 ps=1.966e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m374 222 221 137 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m375 1 19 222 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.764e-11 ad=2.38e-11 ps=7.049e-05 pd=2.97e-05 
+ nrs=0.07 nrd=0.03 
m376 0 214 221 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.806e-11 ad=2.562e-11 ps=2.064e-05 pd=2.29e-05 
+ nrs=0.26 nrd=0.36 
m377 1 214 221 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.211e-11 ad=2.694e-11 ps=3.927e-05 pd=3.57e-05 
+ nrs=0.13 nrd=0.11 
m378 155 223 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.72e-11 ps=1.13e-05 pd=1.966e-05 
+ nrs=0.21 nrd=0.27 
m379 0 167 155 0 nenh l=1.1e-06 w=8e-06 
+ as=1.72e-11 ad=1.32e-11 ps=1.966e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m380 224 223 155 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m381 1 167 224 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.764e-11 ad=2.38e-11 ps=7.049e-05 pd=2.97e-05 
+ nrs=0.07 nrd=0.03 
m382 225 226 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.72e-11 ps=1.13e-05 pd=1.966e-05 
+ nrs=0.21 nrd=0.27 
m383 0 227 225 0 nenh l=1.1e-06 w=8e-06 
+ as=1.72e-11 ad=1.32e-11 ps=1.966e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m384 228 226 225 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m385 1 227 228 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.764e-11 ad=2.38e-11 ps=7.049e-05 pd=2.97e-05 
+ nrs=0.07 nrd=0.03 
m386 0 230 229 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.806e-11 ad=2.562e-11 ps=2.064e-05 pd=2.29e-05 
+ nrs=0.26 nrd=0.36 
m387 1 230 229 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.211e-11 ad=2.694e-11 ps=3.927e-05 pd=3.57e-05 
+ nrs=0.13 nrd=0.11 
m388 231 143 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.72e-11 ps=1.13e-05 pd=1.966e-05 
+ nrs=0.21 nrd=0.27 
m389 0 157 231 0 nenh l=1.1e-06 w=8e-06 
+ as=1.72e-11 ad=1.32e-11 ps=1.966e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m390 232 143 231 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m391 1 157 232 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.764e-11 ad=2.38e-11 ps=7.049e-05 pd=2.97e-05 
+ nrs=0.07 nrd=0.03 
m392 230 173 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.72e-11 ps=1.13e-05 pd=1.966e-05 
+ nrs=0.21 nrd=0.27 
m393 0 143 230 0 nenh l=1.1e-06 w=8e-06 
+ as=1.72e-11 ad=1.32e-11 ps=1.966e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m394 233 173 230 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m395 1 143 233 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.764e-11 ad=2.38e-11 ps=7.049e-05 pd=2.97e-05 
+ nrs=0.07 nrd=0.03 
m396 234 235 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.72e-11 ps=1.13e-05 pd=1.966e-05 
+ nrs=0.21 nrd=0.27 
m397 0 143 234 0 nenh l=1.1e-06 w=8e-06 
+ as=1.72e-11 ad=1.32e-11 ps=1.966e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m398 236 235 234 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m399 1 143 236 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.764e-11 ad=2.38e-11 ps=7.049e-05 pd=2.97e-05 
+ nrs=0.07 nrd=0.03 
m400 0 149 235 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.806e-11 ad=2.562e-11 ps=2.064e-05 pd=2.29e-05 
+ nrs=0.26 nrd=0.36 
m401 1 149 235 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.211e-11 ad=2.694e-11 ps=3.927e-05 pd=3.57e-05 
+ nrs=0.13 nrd=0.11 
m402 237 162 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.72e-11 ps=1.13e-05 pd=1.966e-05 
+ nrs=0.21 nrd=0.27 
m403 0 238 237 0 nenh l=1.1e-06 w=8e-06 
+ as=1.72e-11 ad=1.32e-11 ps=1.966e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m404 239 162 237 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m405 1 238 239 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.764e-11 ad=2.38e-11 ps=7.049e-05 pd=2.97e-05 
+ nrs=0.07 nrd=0.03 
m406 0 237 240 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.806e-11 ad=2.562e-11 ps=2.064e-05 pd=2.29e-05 
+ nrs=0.26 nrd=0.36 
m407 1 237 240 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.211e-11 ad=2.694e-11 ps=3.927e-05 pd=3.57e-05 
+ nrs=0.13 nrd=0.11 
m408 0 242 241 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.806e-11 ad=2.562e-11 ps=2.064e-05 pd=2.29e-05 
+ nrs=0.26 nrd=0.36 
m409 1 242 241 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.211e-11 ad=2.694e-11 ps=3.927e-05 pd=3.57e-05 
+ nrs=0.13 nrd=0.11 
m410 185 241 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.72e-11 ps=1.13e-05 pd=1.966e-05 
+ nrs=0.21 nrd=0.27 
m411 0 162 185 0 nenh l=1.1e-06 w=8e-06 
+ as=1.72e-11 ad=1.32e-11 ps=1.966e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m412 243 241 185 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m413 1 162 243 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.764e-11 ad=2.38e-11 ps=7.049e-05 pd=2.97e-05 
+ nrs=0.07 nrd=0.03 
m414 86 169 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.72e-11 ps=1.13e-05 pd=1.966e-05 
+ nrs=0.21 nrd=0.27 
m415 0 109 86 0 nenh l=1.1e-06 w=8e-06 
+ as=1.72e-11 ad=1.32e-11 ps=1.966e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m416 244 169 86 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m417 1 109 244 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.764e-11 ad=2.38e-11 ps=7.049e-05 pd=2.97e-05 
+ nrs=0.07 nrd=0.03 
m418 245 140 223 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m419 0 139 245 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.44e-11 ad=1.36e-11 ps=3.932e-05 pd=1.77e-05 
+ nrs=0.13 nrd=0.05 
m420 223 140 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.882e-11 ps=1.73e-05 pd=3.524e-05 
+ nrs=0.12 nrd=0.15 
m421 1 139 223 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.882e-11 ad=2.31e-11 ps=3.524e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m422 246 226 247 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m423 0 227 246 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.44e-11 ad=1.36e-11 ps=3.932e-05 pd=1.77e-05 
+ nrs=0.13 nrd=0.05 
m424 247 226 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.882e-11 ps=1.73e-05 pd=3.524e-05 
+ nrs=0.12 nrd=0.15 
m425 1 227 247 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.882e-11 ad=2.31e-11 ps=3.524e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m426 248 229 249 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m427 0 149 248 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.44e-11 ad=1.36e-11 ps=3.932e-05 pd=1.77e-05 
+ nrs=0.13 nrd=0.05 
m428 249 229 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.882e-11 ps=1.73e-05 pd=3.524e-05 
+ nrs=0.12 nrd=0.15 
m429 1 149 249 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.882e-11 ad=2.31e-11 ps=3.524e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m430 0 143 250 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.44e-11 ad=3.008e-11 ps=3.932e-05 pd=3.81e-05 
+ nrs=0.13 nrd=0.12 
m431 251 184 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=3.44e-11 ps=1.77e-05 pd=3.932e-05 
+ nrs=0.05 nrd=0.13 
m432 250 149 251 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.008e-11 ad=1.36e-11 ps=3.81e-05 pd=1.77e-05 
+ nrs=0.12 nrd=0.05 
m433 252 143 250 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=3.5e-11 ps=4.183e-05 pd=6.21e-05 
+ nrs=0.06 nrd=0.04 
m434 1 184 252 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.764e-11 ad=4.62e-11 ps=7.049e-05 pd=4.183e-05 
+ nrs=0.07 nrd=0.06 
m435 252 149 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.764e-11 ps=4.183e-05 pd=7.049e-05 
+ nrs=0.06 nrd=0.07 
m436 253 175 242 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m437 0 238 253 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.44e-11 ad=1.36e-11 ps=3.932e-05 pd=1.77e-05 
+ nrs=0.13 nrd=0.05 
m438 242 175 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.882e-11 ps=1.73e-05 pd=3.524e-05 
+ nrs=0.12 nrd=0.15 
m439 1 238 242 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.882e-11 ad=2.31e-11 ps=3.524e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m440 254 240 182 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m441 0 175 254 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.44e-11 ad=1.36e-11 ps=3.932e-05 pd=1.77e-05 
+ nrs=0.13 nrd=0.05 
m442 182 240 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.882e-11 ps=1.73e-05 pd=3.524e-05 
+ nrs=0.12 nrd=0.15 
m443 1 175 182 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.882e-11 ad=2.31e-11 ps=3.524e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m444 255 257 256 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m445 0 185 255 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.44e-11 ad=2.507e-11 ps=3.932e-05 pd=2.557e-05 
+ nrs=0.13 nrd=0.1 
m446 255 179 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.44e-11 ps=2.557e-05 pd=3.932e-05 
+ nrs=0.1 nrd=0.13 
m447 256 257 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.764e-11 ps=3.13e-05 pd=7.049e-05 
+ nrs=0.06 nrd=0.07 
m448 258 185 256 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m449 1 179 258 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.764e-11 ad=4.62e-11 ps=7.049e-05 pd=3.13e-05 
+ nrs=0.07 nrd=0.06 
m450 259 182 257 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m451 0 179 259 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.44e-11 ad=1.36e-11 ps=3.932e-05 pd=1.77e-05 
+ nrs=0.13 nrd=0.05 
m452 257 182 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.882e-11 ps=1.73e-05 pd=3.524e-05 
+ nrs=0.12 nrd=0.15 
m453 1 179 257 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.882e-11 ad=2.31e-11 ps=3.524e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m454 0 261 260 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.44e-11 ad=3.008e-11 ps=3.932e-05 pd=3.81e-05 
+ nrs=0.13 nrd=0.12 
m455 262 184 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=3.44e-11 ps=1.77e-05 pd=3.932e-05 
+ nrs=0.05 nrd=0.13 
m456 260 234 262 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.008e-11 ad=1.36e-11 ps=3.81e-05 pd=1.77e-05 
+ nrs=0.12 nrd=0.05 
m457 263 261 260 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=3.5e-11 ps=4.183e-05 pd=6.21e-05 
+ nrs=0.06 nrd=0.04 
m458 1 184 263 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.764e-11 ad=4.62e-11 ps=7.049e-05 pd=4.183e-05 
+ nrs=0.07 nrd=0.06 
m459 263 234 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.764e-11 ps=4.183e-05 pd=7.049e-05 
+ nrs=0.06 nrd=0.07 
m460 264 12 265 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m461 0 101 264 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.465e-11 ad=2.507e-11 ps=3.9e-05 pd=2.557e-05 
+ nrs=0.14 nrd=0.1 
m462 264 3 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.465e-11 ps=2.557e-05 pd=3.9e-05 
+ nrs=0.1 nrd=0.14 
m463 265 12 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.755e-11 ps=3.13e-05 pd=7.074e-05 
+ nrs=0.06 nrd=0.07 
m464 266 101 265 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m465 1 3 266 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.755e-11 ad=4.62e-11 ps=7.074e-05 pd=3.13e-05 
+ nrs=0.07 nrd=0.06 
m466 0 265 267 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.819e-11 ad=2.562e-11 ps=2.047e-05 pd=2.29e-05 
+ nrs=0.26 nrd=0.36 
m467 1 265 267 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.206e-11 ad=2.694e-11 ps=3.941e-05 pd=3.57e-05 
+ nrs=0.13 nrd=0.11 
m468 268 270 269 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m469 0 271 268 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.465e-11 ad=2.507e-11 ps=3.9e-05 pd=2.557e-05 
+ nrs=0.14 nrd=0.1 
m470 268 167 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.465e-11 ps=2.557e-05 pd=3.9e-05 
+ nrs=0.1 nrd=0.14 
m471 269 270 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.755e-11 ps=3.13e-05 pd=7.074e-05 
+ nrs=0.06 nrd=0.07 
m472 272 271 269 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m473 1 167 272 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.755e-11 ad=4.62e-11 ps=7.074e-05 pd=3.13e-05 
+ nrs=0.07 nrd=0.06 
m474 273 274 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.732e-11 ps=1.13e-05 pd=1.95e-05 
+ nrs=0.21 nrd=0.27 
m475 0 275 273 0 nenh l=1.1e-06 w=8e-06 
+ as=1.732e-11 ad=1.32e-11 ps=1.95e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m476 276 274 273 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m477 1 275 276 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.755e-11 ad=2.38e-11 ps=7.074e-05 pd=2.97e-05 
+ nrs=0.07 nrd=0.03 
m478 0 273 277 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.819e-11 ad=2.562e-11 ps=2.047e-05 pd=2.29e-05 
+ nrs=0.26 nrd=0.36 
m479 1 273 277 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.206e-11 ad=2.694e-11 ps=3.941e-05 pd=3.57e-05 
+ nrs=0.13 nrd=0.11 
m480 0 277 167 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.819e-11 ad=2.562e-11 ps=2.047e-05 pd=2.29e-05 
+ nrs=0.26 nrd=0.36 
m481 1 277 167 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.206e-11 ad=2.694e-11 ps=3.941e-05 pd=3.57e-05 
+ nrs=0.13 nrd=0.11 
m482 271 113 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.732e-11 ps=1.13e-05 pd=1.95e-05 
+ nrs=0.21 nrd=0.27 
m483 0 109 271 0 nenh l=1.1e-06 w=8e-06 
+ as=1.732e-11 ad=1.32e-11 ps=1.95e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m484 278 113 271 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m485 1 109 278 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.755e-11 ad=2.38e-11 ps=7.074e-05 pd=2.97e-05 
+ nrs=0.07 nrd=0.03 
m486 279 223 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.732e-11 ps=1.13e-05 pd=1.95e-05 
+ nrs=0.21 nrd=0.27 
m487 0 15 279 0 nenh l=1.1e-06 w=8e-06 
+ as=1.732e-11 ad=1.32e-11 ps=1.95e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m488 280 223 279 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m489 1 15 280 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.755e-11 ad=2.38e-11 ps=7.074e-05 pd=2.97e-05 
+ nrs=0.07 nrd=0.03 
m490 281 282 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.732e-11 ps=1.13e-05 pd=1.95e-05 
+ nrs=0.21 nrd=0.27 
m491 0 283 281 0 nenh l=1.1e-06 w=8e-06 
+ as=1.732e-11 ad=1.32e-11 ps=1.95e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m492 284 282 281 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m493 1 283 284 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.755e-11 ad=2.38e-11 ps=7.074e-05 pd=2.97e-05 
+ nrs=0.07 nrd=0.03 
m494 0 124 285 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.819e-11 ad=2.562e-11 ps=2.047e-05 pd=2.29e-05 
+ nrs=0.26 nrd=0.36 
m495 1 124 285 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.206e-11 ad=2.694e-11 ps=3.941e-05 pd=3.57e-05 
+ nrs=0.13 nrd=0.11 
m496 286 287 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.732e-11 ps=1.13e-05 pd=1.95e-05 
+ nrs=0.21 nrd=0.27 
m497 0 288 286 0 nenh l=1.1e-06 w=8e-06 
+ as=1.732e-11 ad=1.32e-11 ps=1.95e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m498 289 287 286 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m499 1 288 289 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.755e-11 ad=2.38e-11 ps=7.074e-05 pd=2.97e-05 
+ nrs=0.07 nrd=0.03 
m500 290 291 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.732e-11 ps=1.13e-05 pd=1.95e-05 
+ nrs=0.21 nrd=0.27 
m501 0 288 290 0 nenh l=1.1e-06 w=8e-06 
+ as=1.732e-11 ad=1.32e-11 ps=1.95e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m502 292 291 290 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m503 1 288 292 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.755e-11 ad=2.38e-11 ps=7.074e-05 pd=2.97e-05 
+ nrs=0.07 nrd=0.03 
m504 0 293 291 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.819e-11 ad=2.562e-11 ps=2.047e-05 pd=2.29e-05 
+ nrs=0.26 nrd=0.36 
m505 1 293 291 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.206e-11 ad=2.694e-11 ps=3.941e-05 pd=3.57e-05 
+ nrs=0.13 nrd=0.11 
m506 288 294 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.732e-11 ps=1.13e-05 pd=1.95e-05 
+ nrs=0.21 nrd=0.27 
m507 0 295 288 0 nenh l=1.1e-06 w=8e-06 
+ as=1.732e-11 ad=1.32e-11 ps=1.95e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m508 296 294 288 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m509 1 295 296 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.755e-11 ad=2.38e-11 ps=7.074e-05 pd=2.97e-05 
+ nrs=0.07 nrd=0.03 
m510 0 286 297 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.819e-11 ad=2.562e-11 ps=2.047e-05 pd=2.29e-05 
+ nrs=0.26 nrd=0.36 
m511 1 286 297 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.206e-11 ad=2.694e-11 ps=3.941e-05 pd=3.57e-05 
+ nrs=0.13 nrd=0.11 
m512 298 299 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.732e-11 ps=1.13e-05 pd=1.95e-05 
+ nrs=0.21 nrd=0.27 
m513 0 300 298 0 nenh l=1.1e-06 w=8e-06 
+ as=1.732e-11 ad=1.32e-11 ps=1.95e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m514 301 299 298 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m515 1 300 301 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.755e-11 ad=2.38e-11 ps=7.074e-05 pd=2.97e-05 
+ nrs=0.07 nrd=0.03 
m516 0 303 302 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.819e-11 ad=2.562e-11 ps=2.047e-05 pd=2.29e-05 
+ nrs=0.26 nrd=0.36 
m517 1 303 302 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.206e-11 ad=2.694e-11 ps=3.941e-05 pd=3.57e-05 
+ nrs=0.13 nrd=0.11 
m518 304 249 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.732e-11 ps=1.13e-05 pd=1.95e-05 
+ nrs=0.21 nrd=0.27 
m519 0 302 304 0 nenh l=1.1e-06 w=8e-06 
+ as=1.732e-11 ad=1.32e-11 ps=1.95e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m520 305 249 304 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m521 1 302 305 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.755e-11 ad=2.38e-11 ps=7.074e-05 pd=2.97e-05 
+ nrs=0.07 nrd=0.03 
m522 306 307 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.732e-11 ps=1.13e-05 pd=1.95e-05 
+ nrs=0.21 nrd=0.27 
m523 0 225 306 0 nenh l=1.1e-06 w=8e-06 
+ as=1.732e-11 ad=1.32e-11 ps=1.95e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m524 308 307 306 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m525 1 225 308 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.755e-11 ad=2.38e-11 ps=7.074e-05 pd=2.97e-05 
+ nrs=0.07 nrd=0.03 
m526 0 175 309 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.819e-11 ad=2.562e-11 ps=2.047e-05 pd=2.29e-05 
+ nrs=0.26 nrd=0.36 
m527 1 175 309 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.206e-11 ad=2.694e-11 ps=3.941e-05 pd=3.57e-05 
+ nrs=0.13 nrd=0.11 
m528 0 162 310 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.819e-11 ad=2.562e-11 ps=2.047e-05 pd=2.29e-05 
+ nrs=0.26 nrd=0.36 
m529 1 162 310 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.206e-11 ad=2.694e-11 ps=3.941e-05 pd=3.57e-05 
+ nrs=0.13 nrd=0.11 
m530 311 309 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.732e-11 ps=1.13e-05 pd=1.95e-05 
+ nrs=0.21 nrd=0.27 
m531 0 162 311 0 nenh l=1.1e-06 w=8e-06 
+ as=1.732e-11 ad=1.32e-11 ps=1.95e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m532 312 309 311 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m533 1 162 312 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.755e-11 ad=2.38e-11 ps=7.074e-05 pd=2.97e-05 
+ nrs=0.07 nrd=0.03 
m534 313 307 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.732e-11 ps=1.13e-05 pd=1.95e-05 
+ nrs=0.21 nrd=0.27 
m535 0 238 313 0 nenh l=1.1e-06 w=8e-06 
+ as=1.732e-11 ad=1.32e-11 ps=1.95e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m536 314 307 313 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m537 1 238 314 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.755e-11 ad=2.38e-11 ps=7.074e-05 pd=2.97e-05 
+ nrs=0.07 nrd=0.03 
m538 0 83 315 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.819e-11 ad=2.562e-11 ps=2.047e-05 pd=2.29e-05 
+ nrs=0.26 nrd=0.36 
m539 1 83 315 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.206e-11 ad=2.694e-11 ps=3.941e-05 pd=3.57e-05 
+ nrs=0.13 nrd=0.11 
m540 316 315 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.732e-11 ps=1.13e-05 pd=1.95e-05 
+ nrs=0.21 nrd=0.27 
m541 0 70 316 0 nenh l=1.1e-06 w=8e-06 
+ as=1.732e-11 ad=1.32e-11 ps=1.95e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m542 317 315 316 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m543 1 70 317 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.755e-11 ad=2.38e-11 ps=7.074e-05 pd=2.97e-05 
+ nrs=0.07 nrd=0.03 
m544 318 319 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.732e-11 ps=1.13e-05 pd=1.95e-05 
+ nrs=0.21 nrd=0.27 
m545 0 320 318 0 nenh l=1.1e-06 w=8e-06 
+ as=1.732e-11 ad=1.32e-11 ps=1.95e-05 pd=1.13e-05 
+ nrs=0.27 nrd=0.21 
m546 321 319 318 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m547 1 320 321 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.755e-11 ad=2.38e-11 ps=7.074e-05 pd=2.97e-05 
+ nrs=0.07 nrd=0.03 
m548 322 271 270 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m549 0 167 322 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.465e-11 ad=1.36e-11 ps=3.9e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m550 270 271 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.878e-11 ps=1.73e-05 pd=3.537e-05 
+ nrs=0.12 nrd=0.15 
m551 1 167 270 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.878e-11 ad=2.31e-11 ps=3.537e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m552 323 275 324 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m553 0 279 323 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.465e-11 ad=1.36e-11 ps=3.9e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m554 324 275 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.878e-11 ps=1.73e-05 pd=3.537e-05 
+ nrs=0.12 nrd=0.15 
m555 1 279 324 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.878e-11 ad=2.31e-11 ps=3.537e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m556 325 274 326 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m557 0 279 325 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.465e-11 ad=1.36e-11 ps=3.9e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m558 326 274 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.878e-11 ps=1.73e-05 pd=3.537e-05 
+ nrs=0.12 nrd=0.15 
m559 1 279 326 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.878e-11 ad=2.31e-11 ps=3.537e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m560 327 282 287 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m561 0 283 327 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.465e-11 ad=1.36e-11 ps=3.9e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m562 287 282 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.878e-11 ps=1.73e-05 pd=3.537e-05 
+ nrs=0.12 nrd=0.15 
m563 1 283 287 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.878e-11 ad=2.31e-11 ps=3.537e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m564 328 294 293 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m565 0 295 328 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.465e-11 ad=1.36e-11 ps=3.9e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m566 293 294 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.878e-11 ps=1.73e-05 pd=3.537e-05 
+ nrs=0.12 nrd=0.15 
m567 1 295 293 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.878e-11 ad=2.31e-11 ps=3.537e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m568 329 297 330 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m569 0 293 329 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.465e-11 ad=1.36e-11 ps=3.9e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m570 330 297 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.878e-11 ps=1.73e-05 pd=3.537e-05 
+ nrs=0.12 nrd=0.15 
m571 1 293 330 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.878e-11 ad=2.31e-11 ps=3.537e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m572 331 299 332 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m573 0 300 331 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.465e-11 ad=1.36e-11 ps=3.9e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m574 332 299 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.878e-11 ps=1.73e-05 pd=3.537e-05 
+ nrs=0.12 nrd=0.15 
m575 1 300 332 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.878e-11 ad=2.31e-11 ps=3.537e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m576 333 231 303 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m577 0 309 333 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.465e-11 ad=1.36e-11 ps=3.9e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m578 303 231 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.878e-11 ps=1.73e-05 pd=3.537e-05 
+ nrs=0.12 nrd=0.15 
m579 1 309 303 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.878e-11 ad=2.31e-11 ps=3.537e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m580 334 231 307 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m581 0 310 334 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.465e-11 ad=1.36e-11 ps=3.9e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m582 307 231 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.878e-11 ps=1.73e-05 pd=3.537e-05 
+ nrs=0.12 nrd=0.15 
m583 1 310 307 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.878e-11 ad=2.31e-11 ps=3.537e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m584 335 319 336 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m585 0 320 335 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.465e-11 ad=1.36e-11 ps=3.9e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m586 336 319 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.878e-11 ps=1.73e-05 pd=3.537e-05 
+ nrs=0.12 nrd=0.15 
m587 1 320 336 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.878e-11 ad=2.31e-11 ps=3.537e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m588 0 318 337 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.465e-11 ad=3.008e-11 ps=3.9e-05 pd=3.81e-05 
+ nrs=0.14 nrd=0.12 
m589 338 339 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=3.465e-11 ps=1.77e-05 pd=3.9e-05 
+ nrs=0.05 nrd=0.14 
m590 337 336 338 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.008e-11 ad=1.36e-11 ps=3.81e-05 pd=1.77e-05 
+ nrs=0.12 nrd=0.05 
m591 340 318 337 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=3.5e-11 ps=4.183e-05 pd=6.21e-05 
+ nrs=0.06 nrd=0.04 
m592 1 339 340 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.755e-11 ad=4.62e-11 ps=7.074e-05 pd=4.183e-05 
+ nrs=0.07 nrd=0.06 
m593 340 336 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.755e-11 ps=4.183e-05 pd=7.074e-05 
+ nrs=0.06 nrd=0.07 
m594 341 343 342 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m595 0 337 341 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.465e-11 ad=2.507e-11 ps=3.9e-05 pd=2.557e-05 
+ nrs=0.14 nrd=0.1 
m596 341 344 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.465e-11 ps=2.557e-05 pd=3.9e-05 
+ nrs=0.1 nrd=0.14 
m597 342 343 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.755e-11 ps=3.13e-05 pd=7.074e-05 
+ nrs=0.06 nrd=0.07 
m598 345 337 342 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m599 1 344 345 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.755e-11 ad=4.62e-11 ps=7.074e-05 pd=3.13e-05 
+ nrs=0.07 nrd=0.06 
m600 346 344 343 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m601 0 347 346 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.465e-11 ad=2.507e-11 ps=3.9e-05 pd=2.557e-05 
+ nrs=0.14 nrd=0.1 
m602 346 348 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.465e-11 ps=2.557e-05 pd=3.9e-05 
+ nrs=0.1 nrd=0.14 
m603 343 344 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.755e-11 ps=3.13e-05 pd=7.074e-05 
+ nrs=0.06 nrd=0.07 
m604 349 347 343 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m605 1 348 349 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.755e-11 ad=4.62e-11 ps=7.074e-05 pd=3.13e-05 
+ nrs=0.07 nrd=0.06 
m606 350 351 344 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m607 0 352 350 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.465e-11 ad=2.507e-11 ps=3.9e-05 pd=2.557e-05 
+ nrs=0.14 nrd=0.1 
m608 350 353 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.465e-11 ps=2.557e-05 pd=3.9e-05 
+ nrs=0.1 nrd=0.14 
m609 344 351 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.755e-11 ps=3.13e-05 pd=7.074e-05 
+ nrs=0.06 nrd=0.07 
m610 354 352 344 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m611 1 353 354 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.755e-11 ad=4.62e-11 ps=7.074e-05 pd=3.13e-05 
+ nrs=0.07 nrd=0.06 
m612 355 352 351 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m613 0 353 355 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.465e-11 ad=1.36e-11 ps=3.9e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m614 351 352 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.878e-11 ps=1.73e-05 pd=3.537e-05 
+ nrs=0.12 nrd=0.15 
m615 1 353 351 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.878e-11 ad=2.31e-11 ps=3.537e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m616 356 358 357 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m617 0 86 356 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.465e-11 ad=2.507e-11 ps=3.9e-05 pd=2.557e-05 
+ nrs=0.14 nrd=0.1 
m618 356 100 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.465e-11 ps=2.557e-05 pd=3.9e-05 
+ nrs=0.1 nrd=0.14 
m619 357 358 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.755e-11 ps=3.13e-05 pd=7.074e-05 
+ nrs=0.06 nrd=0.07 
m620 359 86 357 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m621 1 100 359 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.755e-11 ad=4.62e-11 ps=7.074e-05 pd=3.13e-05 
+ nrs=0.07 nrd=0.06 
m622 0 173 186 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.819e-11 ad=2.562e-11 ps=2.047e-05 pd=2.29e-05 
+ nrs=0.26 nrd=0.36 
m623 1 173 186 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.206e-11 ad=2.694e-11 ps=3.941e-05 pd=3.57e-05 
+ nrs=0.13 nrd=0.11 
m624 0 234 261 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.465e-11 ad=3.008e-11 ps=3.9e-05 pd=3.81e-05 
+ nrs=0.14 nrd=0.12 
m625 360 181 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=3.465e-11 ps=1.77e-05 pd=3.9e-05 
+ nrs=0.05 nrd=0.14 
m626 261 173 360 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.008e-11 ad=1.36e-11 ps=3.81e-05 pd=1.77e-05 
+ nrs=0.12 nrd=0.05 
m627 361 234 261 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=3.5e-11 ps=4.183e-05 pd=6.21e-05 
+ nrs=0.06 nrd=0.04 
m628 1 181 361 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.755e-11 ad=4.62e-11 ps=7.074e-05 pd=4.183e-05 
+ nrs=0.07 nrd=0.06 
m629 361 173 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.755e-11 ps=4.183e-05 pd=7.074e-05 
+ nrs=0.06 nrd=0.07 
m630 362 363 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.821e-11 ps=1.13e-05 pd=1.961e-05 
+ nrs=0.21 nrd=0.28 
m631 0 364 362 0 nenh l=1.1e-06 w=8e-06 
+ as=1.821e-11 ad=1.32e-11 ps=1.961e-05 pd=1.13e-05 
+ nrs=0.28 nrd=0.21 
m632 365 363 362 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m633 1 364 365 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.08e-11 ad=2.38e-11 ps=7.147e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m634 0 362 366 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.912e-11 ad=2.562e-11 ps=2.059e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m635 1 362 366 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.387e-11 ad=2.694e-11 ps=3.982e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m636 0 366 274 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.642e-11 ad=3.008e-11 ps=3.922e-05 pd=3.81e-05 
+ nrs=0.14 nrd=0.12 
m637 367 192 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=3.642e-11 ps=1.77e-05 pd=3.922e-05 
+ nrs=0.05 nrd=0.14 
m638 274 267 367 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.008e-11 ad=1.36e-11 ps=3.81e-05 pd=1.77e-05 
+ nrs=0.12 nrd=0.05 
m639 368 366 274 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=3.5e-11 ps=4.183e-05 pd=6.21e-05 
+ nrs=0.06 nrd=0.04 
m640 1 192 368 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.08e-11 ad=4.62e-11 ps=7.147e-05 pd=4.183e-05 
+ nrs=0.08 nrd=0.06 
m641 368 267 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=6.08e-11 ps=4.183e-05 pd=7.147e-05 
+ nrs=0.06 nrd=0.08 
m642 0 370 369 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.912e-11 ad=2.562e-11 ps=2.059e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m643 1 370 369 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.387e-11 ad=2.694e-11 ps=3.982e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m644 0 372 371 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.912e-11 ad=2.562e-11 ps=2.059e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m645 1 372 371 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.387e-11 ad=2.694e-11 ps=3.982e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m646 373 330 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.821e-11 ps=1.13e-05 pd=1.961e-05 
+ nrs=0.21 nrd=0.28 
m647 0 371 373 0 nenh l=1.1e-06 w=8e-06 
+ as=1.821e-11 ad=1.32e-11 ps=1.961e-05 pd=1.13e-05 
+ nrs=0.28 nrd=0.21 
m648 374 330 373 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m649 1 371 374 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.08e-11 ad=2.38e-11 ps=7.147e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m650 375 267 370 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m651 0 192 375 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.642e-11 ad=1.36e-11 ps=3.922e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m652 370 267 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=3.04e-11 ps=1.73e-05 pd=3.574e-05 
+ nrs=0.12 nrd=0.16 
m653 1 192 370 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.04e-11 ad=2.31e-11 ps=3.574e-05 pd=1.73e-05 
+ nrs=0.16 nrd=0.12 
m654 376 377 372 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m655 0 378 376 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.642e-11 ad=1.36e-11 ps=3.922e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m656 372 377 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=3.04e-11 ps=1.73e-05 pd=3.574e-05 
+ nrs=0.12 nrd=0.16 
m657 1 378 372 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.04e-11 ad=2.31e-11 ps=3.574e-05 pd=1.73e-05 
+ nrs=0.16 nrd=0.12 
m658 377 288 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.821e-11 ps=1.13e-05 pd=1.961e-05 
+ nrs=0.21 nrd=0.28 
m659 0 281 377 0 nenh l=1.1e-06 w=8e-06 
+ as=1.821e-11 ad=1.32e-11 ps=1.961e-05 pd=1.13e-05 
+ nrs=0.28 nrd=0.21 
m660 379 288 377 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m661 1 281 379 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.08e-11 ad=2.38e-11 ps=7.147e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m662 0 298 380 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.912e-11 ad=2.562e-11 ps=2.059e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m663 1 298 380 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.387e-11 ad=2.694e-11 ps=3.982e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m664 0 281 381 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.912e-11 ad=2.562e-11 ps=2.059e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m665 1 281 381 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.387e-11 ad=2.694e-11 ps=3.982e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m666 382 377 363 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m667 0 380 382 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.642e-11 ad=1.36e-11 ps=3.922e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m668 363 377 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=3.04e-11 ps=1.73e-05 pd=3.574e-05 
+ nrs=0.12 nrd=0.16 
m669 1 380 363 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.04e-11 ad=2.31e-11 ps=3.574e-05 pd=1.73e-05 
+ nrs=0.16 nrd=0.12 
m670 383 287 384 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m671 0 381 383 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.642e-11 ad=1.36e-11 ps=3.922e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m672 384 287 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=3.04e-11 ps=1.73e-05 pd=3.574e-05 
+ nrs=0.12 nrd=0.16 
m673 1 381 384 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.04e-11 ad=2.31e-11 ps=3.574e-05 pd=1.73e-05 
+ nrs=0.16 nrd=0.12 
m674 0 287 385 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.912e-11 ad=2.562e-11 ps=2.059e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m675 1 287 385 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.387e-11 ad=2.694e-11 ps=3.982e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m676 386 387 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.821e-11 ps=1.13e-05 pd=1.961e-05 
+ nrs=0.21 nrd=0.28 
m677 0 298 386 0 nenh l=1.1e-06 w=8e-06 
+ as=1.821e-11 ad=1.32e-11 ps=1.961e-05 pd=1.13e-05 
+ nrs=0.28 nrd=0.21 
m678 388 387 386 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m679 1 298 388 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.08e-11 ad=2.38e-11 ps=7.147e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m680 0 389 387 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.912e-11 ad=2.562e-11 ps=2.059e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m681 1 389 387 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.387e-11 ad=2.694e-11 ps=3.982e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m682 390 298 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.821e-11 ps=1.13e-05 pd=1.961e-05 
+ nrs=0.21 nrd=0.28 
m683 0 369 390 0 nenh l=1.1e-06 w=8e-06 
+ as=1.821e-11 ad=1.32e-11 ps=1.961e-05 pd=1.13e-05 
+ nrs=0.28 nrd=0.21 
m684 391 298 390 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m685 1 369 391 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.08e-11 ad=2.38e-11 ps=7.147e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m686 0 332 378 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.912e-11 ad=2.562e-11 ps=2.059e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m687 1 332 378 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.387e-11 ad=2.694e-11 ps=3.982e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m688 392 378 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.821e-11 ps=1.13e-05 pd=1.961e-05 
+ nrs=0.21 nrd=0.28 
m689 0 298 392 0 nenh l=1.1e-06 w=8e-06 
+ as=1.821e-11 ad=1.32e-11 ps=1.961e-05 pd=1.13e-05 
+ nrs=0.28 nrd=0.21 
m690 393 378 392 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m691 1 298 393 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.08e-11 ad=2.38e-11 ps=7.147e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m692 0 57 394 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.912e-11 ad=2.562e-11 ps=2.059e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m693 1 57 394 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.387e-11 ad=2.694e-11 ps=3.982e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m694 0 288 395 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.642e-11 ad=3.008e-11 ps=3.922e-05 pd=3.81e-05 
+ nrs=0.14 nrd=0.12 
m695 396 397 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=3.642e-11 ps=1.77e-05 pd=3.922e-05 
+ nrs=0.05 nrd=0.14 
m696 395 293 396 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.008e-11 ad=1.36e-11 ps=3.81e-05 pd=1.77e-05 
+ nrs=0.12 nrd=0.05 
m697 398 288 395 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=3.5e-11 ps=4.183e-05 pd=6.21e-05 
+ nrs=0.06 nrd=0.04 
m698 1 397 398 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.08e-11 ad=4.62e-11 ps=7.147e-05 pd=4.183e-05 
+ nrs=0.08 nrd=0.06 
m699 398 293 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=6.08e-11 ps=4.183e-05 pd=7.147e-05 
+ nrs=0.06 nrd=0.08 
m700 399 381 397 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m701 0 386 399 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.642e-11 ad=2.507e-11 ps=3.922e-05 pd=2.557e-05 
+ nrs=0.14 nrd=0.1 
m702 399 385 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.642e-11 ps=2.557e-05 pd=3.922e-05 
+ nrs=0.1 nrd=0.14 
m703 397 381 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=6.08e-11 ps=3.13e-05 pd=7.147e-05 
+ nrs=0.06 nrd=0.08 
m704 400 386 397 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m705 1 385 400 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.08e-11 ad=4.62e-11 ps=7.147e-05 pd=3.13e-05 
+ nrs=0.08 nrd=0.06 
m706 401 332 389 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m707 0 369 401 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.642e-11 ad=1.36e-11 ps=3.922e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m708 389 332 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=3.04e-11 ps=1.73e-05 pd=3.574e-05 
+ nrs=0.12 nrd=0.16 
m709 1 369 389 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.04e-11 ad=2.31e-11 ps=3.574e-05 pd=1.73e-05 
+ nrs=0.16 nrd=0.12 
m710 402 324 403 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m711 0 394 402 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.642e-11 ad=1.36e-11 ps=3.922e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m712 403 324 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=3.04e-11 ps=1.73e-05 pd=3.574e-05 
+ nrs=0.12 nrd=0.16 
m713 1 394 403 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.04e-11 ad=2.31e-11 ps=3.574e-05 pd=1.73e-05 
+ nrs=0.16 nrd=0.12 
m714 0 405 404 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.912e-11 ad=2.562e-11 ps=2.059e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m715 1 405 404 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.387e-11 ad=2.694e-11 ps=3.982e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m716 0 406 238 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.912e-11 ad=2.562e-11 ps=2.059e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m717 1 406 238 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.387e-11 ad=2.694e-11 ps=3.982e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m718 0 225 407 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.912e-11 ad=2.562e-11 ps=2.059e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m719 1 225 407 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.387e-11 ad=2.694e-11 ps=3.982e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m720 0 304 408 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.912e-11 ad=2.562e-11 ps=2.059e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m721 1 304 408 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.387e-11 ad=2.694e-11 ps=3.982e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m722 0 336 348 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.912e-11 ad=2.562e-11 ps=2.059e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m723 1 336 348 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.387e-11 ad=2.694e-11 ps=3.982e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m724 409 348 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.821e-11 ps=1.13e-05 pd=1.961e-05 
+ nrs=0.21 nrd=0.28 
m725 0 318 409 0 nenh l=1.1e-06 w=8e-06 
+ as=1.821e-11 ad=1.32e-11 ps=1.961e-05 pd=1.13e-05 
+ nrs=0.28 nrd=0.21 
m726 410 348 409 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m727 1 318 410 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.08e-11 ad=2.38e-11 ps=7.147e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m728 347 411 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.821e-11 ps=1.13e-05 pd=1.961e-05 
+ nrs=0.21 nrd=0.28 
m729 0 318 347 0 nenh l=1.1e-06 w=8e-06 
+ as=1.821e-11 ad=1.32e-11 ps=1.961e-05 pd=1.13e-05 
+ nrs=0.28 nrd=0.21 
m730 412 411 347 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m731 1 318 412 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.08e-11 ad=2.38e-11 ps=7.147e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m732 0 414 413 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.912e-11 ad=2.562e-11 ps=2.059e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m733 1 414 413 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.387e-11 ad=2.694e-11 ps=3.982e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m734 0 416 415 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.912e-11 ad=2.562e-11 ps=2.059e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m735 1 416 415 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.387e-11 ad=2.694e-11 ps=3.982e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m736 414 417 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.821e-11 ps=1.13e-05 pd=1.961e-05 
+ nrs=0.21 nrd=0.28 
m737 0 418 414 0 nenh l=1.1e-06 w=8e-06 
+ as=1.821e-11 ad=1.32e-11 ps=1.961e-05 pd=1.13e-05 
+ nrs=0.28 nrd=0.21 
m738 419 417 414 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m739 1 418 419 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.08e-11 ad=2.38e-11 ps=7.147e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m740 0 260 420 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.912e-11 ad=2.562e-11 ps=2.059e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m741 1 260 420 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.387e-11 ad=2.694e-11 ps=3.982e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m742 421 324 405 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m743 0 394 421 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.642e-11 ad=1.36e-11 ps=3.922e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m744 405 324 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=3.04e-11 ps=1.73e-05 pd=3.574e-05 
+ nrs=0.12 nrd=0.16 
m745 1 394 405 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.04e-11 ad=2.31e-11 ps=3.574e-05 pd=1.73e-05 
+ nrs=0.16 nrd=0.12 
m746 422 326 406 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m747 0 404 422 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.642e-11 ad=1.36e-11 ps=3.922e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m748 406 326 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=3.04e-11 ps=1.73e-05 pd=3.574e-05 
+ nrs=0.12 nrd=0.16 
m749 1 404 406 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.04e-11 ad=2.31e-11 ps=3.574e-05 pd=1.73e-05 
+ nrs=0.16 nrd=0.12 
m750 423 247 424 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m751 0 304 423 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.642e-11 ad=2.507e-11 ps=3.922e-05 pd=2.557e-05 
+ nrs=0.14 nrd=0.1 
m752 423 225 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.642e-11 ps=2.557e-05 pd=3.922e-05 
+ nrs=0.1 nrd=0.14 
m753 424 247 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=6.08e-11 ps=3.13e-05 pd=7.147e-05 
+ nrs=0.06 nrd=0.08 
m754 425 304 424 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m755 1 225 425 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.08e-11 ad=4.62e-11 ps=7.147e-05 pd=3.13e-05 
+ nrs=0.08 nrd=0.06 
m756 426 247 427 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m757 0 407 426 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.642e-11 ad=1.36e-11 ps=3.922e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m758 427 247 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=3.04e-11 ps=1.73e-05 pd=3.574e-05 
+ nrs=0.12 nrd=0.16 
m759 1 407 427 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.04e-11 ad=2.31e-11 ps=3.574e-05 pd=1.73e-05 
+ nrs=0.16 nrd=0.12 
m760 428 427 429 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m761 0 313 428 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.642e-11 ad=2.507e-11 ps=3.922e-05 pd=2.557e-05 
+ nrs=0.14 nrd=0.1 
m762 428 408 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.642e-11 ps=2.557e-05 pd=3.922e-05 
+ nrs=0.1 nrd=0.14 
m763 429 427 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=6.08e-11 ps=3.13e-05 pd=7.147e-05 
+ nrs=0.06 nrd=0.08 
m764 430 313 429 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m765 1 408 430 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.08e-11 ad=4.62e-11 ps=7.147e-05 pd=3.13e-05 
+ nrs=0.08 nrd=0.06 
m766 431 429 432 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m767 0 250 431 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.642e-11 ad=2.507e-11 ps=3.922e-05 pd=2.557e-05 
+ nrs=0.14 nrd=0.1 
m768 431 427 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.642e-11 ps=2.557e-05 pd=3.922e-05 
+ nrs=0.1 nrd=0.14 
m769 432 429 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=6.08e-11 ps=3.13e-05 pd=7.147e-05 
+ nrs=0.06 nrd=0.08 
m770 433 250 432 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m771 1 427 433 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.08e-11 ad=4.62e-11 ps=7.147e-05 pd=3.13e-05 
+ nrs=0.08 nrd=0.06 
m772 434 339 435 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m773 0 409 434 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.642e-11 ad=1.36e-11 ps=3.922e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m774 435 339 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=3.04e-11 ps=1.73e-05 pd=3.574e-05 
+ nrs=0.12 nrd=0.16 
m775 1 409 435 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.04e-11 ad=2.31e-11 ps=3.574e-05 pd=1.73e-05 
+ nrs=0.16 nrd=0.12 
m776 436 435 437 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m777 0 411 436 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.642e-11 ad=2.507e-11 ps=3.922e-05 pd=2.557e-05 
+ nrs=0.14 nrd=0.1 
m778 436 409 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.642e-11 ps=2.557e-05 pd=3.922e-05 
+ nrs=0.1 nrd=0.14 
m779 437 435 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=6.08e-11 ps=3.13e-05 pd=7.147e-05 
+ nrs=0.06 nrd=0.08 
m780 438 411 437 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m781 1 409 438 1 penh l=1.1e-06 w=2.8e-05 
+ as=6.08e-11 ad=4.62e-11 ps=7.147e-05 pd=3.13e-05 
+ nrs=0.08 nrd=0.06 
m782 439 417 416 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m783 0 418 439 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.642e-11 ad=1.36e-11 ps=3.922e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m784 416 417 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=3.04e-11 ps=1.73e-05 pd=3.574e-05 
+ nrs=0.12 nrd=0.16 
m785 1 418 416 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.04e-11 ad=2.31e-11 ps=3.574e-05 pd=1.73e-05 
+ nrs=0.16 nrd=0.12 
m786 364 440 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.804e-11 ps=1.13e-05 pd=1.788e-05 
+ nrs=0.21 nrd=0.28 
m787 0 441 364 0 nenh l=1.1e-06 w=8e-06 
+ as=1.804e-11 ad=1.32e-11 ps=1.788e-05 pd=1.13e-05 
+ nrs=0.28 nrd=0.21 
m788 442 440 364 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m789 1 441 442 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.938e-11 ad=2.38e-11 ps=6.998e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m790 0 364 443 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.895e-11 ad=2.562e-11 ps=1.878e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m791 1 364 443 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.308e-11 ad=2.694e-11 ps=3.899e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m792 444 440 445 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m793 0 441 444 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.609e-11 ad=1.36e-11 ps=3.577e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m794 445 440 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.969e-11 ps=1.73e-05 pd=3.499e-05 
+ nrs=0.12 nrd=0.15 
m795 1 441 445 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.969e-11 ad=2.31e-11 ps=3.499e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m796 446 445 447 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m797 0 443 446 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.609e-11 ad=1.36e-11 ps=3.577e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m798 447 445 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.969e-11 ps=1.73e-05 pd=3.499e-05 
+ nrs=0.12 nrd=0.15 
m799 1 443 447 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.969e-11 ad=2.31e-11 ps=3.499e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m800 448 450 449 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m801 0 395 448 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.609e-11 ad=2.507e-11 ps=3.577e-05 pd=2.557e-05 
+ nrs=0.14 nrd=0.1 
m802 448 447 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.609e-11 ps=2.557e-05 pd=3.577e-05 
+ nrs=0.1 nrd=0.14 
m803 449 450 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.938e-11 ps=3.13e-05 pd=6.998e-05 
+ nrs=0.06 nrd=0.08 
m804 451 395 449 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m805 1 447 451 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.938e-11 ad=4.62e-11 ps=6.998e-05 pd=3.13e-05 
+ nrs=0.08 nrd=0.06 
m806 452 445 275 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m807 0 373 452 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.609e-11 ad=2.507e-11 ps=3.577e-05 pd=2.557e-05 
+ nrs=0.14 nrd=0.1 
m808 452 364 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.609e-11 ps=2.557e-05 pd=3.577e-05 
+ nrs=0.1 nrd=0.14 
m809 275 445 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.938e-11 ps=3.13e-05 pd=6.998e-05 
+ nrs=0.06 nrd=0.08 
m810 453 373 275 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m811 1 364 453 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.938e-11 ad=4.62e-11 ps=6.998e-05 pd=3.13e-05 
+ nrs=0.08 nrd=0.06 
m812 0 373 454 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.895e-11 ad=2.562e-11 ps=1.878e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m813 1 373 454 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.308e-11 ad=2.694e-11 ps=3.899e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m814 455 363 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.804e-11 ps=1.13e-05 pd=1.788e-05 
+ nrs=0.21 nrd=0.28 
m815 0 369 455 0 nenh l=1.1e-06 w=8e-06 
+ as=1.804e-11 ad=1.32e-11 ps=1.788e-05 pd=1.13e-05 
+ nrs=0.28 nrd=0.21 
m816 456 363 455 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m817 1 369 456 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.938e-11 ad=2.38e-11 ps=6.998e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m818 457 459 458 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m819 0 386 457 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.609e-11 ad=2.507e-11 ps=3.577e-05 pd=2.557e-05 
+ nrs=0.14 nrd=0.1 
m820 457 384 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.609e-11 ps=2.557e-05 pd=3.577e-05 
+ nrs=0.1 nrd=0.14 
m821 458 459 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.938e-11 ps=3.13e-05 pd=6.998e-05 
+ nrs=0.06 nrd=0.08 
m822 460 386 458 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m823 1 384 460 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.938e-11 ad=4.62e-11 ps=6.998e-05 pd=3.13e-05 
+ nrs=0.08 nrd=0.06 
m824 461 447 450 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m825 0 455 461 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.609e-11 ad=2.507e-11 ps=3.577e-05 pd=2.557e-05 
+ nrs=0.14 nrd=0.1 
m826 461 454 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.609e-11 ps=2.557e-05 pd=3.577e-05 
+ nrs=0.1 nrd=0.14 
m827 450 447 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.938e-11 ps=3.13e-05 pd=6.998e-05 
+ nrs=0.06 nrd=0.08 
m828 462 455 450 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m829 1 454 462 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.938e-11 ad=4.62e-11 ps=6.998e-05 pd=3.13e-05 
+ nrs=0.08 nrd=0.06 
m830 463 464 459 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m831 0 384 463 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.609e-11 ad=1.36e-11 ps=3.577e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m832 459 464 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.969e-11 ps=1.73e-05 pd=3.499e-05 
+ nrs=0.12 nrd=0.15 
m833 1 384 459 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.969e-11 ad=2.31e-11 ps=3.499e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m834 465 464 466 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m835 0 381 465 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.609e-11 ad=1.36e-11 ps=3.577e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m836 466 464 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.969e-11 ps=1.73e-05 pd=3.499e-05 
+ nrs=0.12 nrd=0.15 
m837 1 381 466 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.969e-11 ad=2.31e-11 ps=3.499e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m838 0 468 467 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.895e-11 ad=2.562e-11 ps=1.878e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m839 1 468 467 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.308e-11 ad=2.694e-11 ps=3.899e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m840 0 290 469 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.609e-11 ad=3.008e-11 ps=3.577e-05 pd=3.81e-05 
+ nrs=0.14 nrd=0.12 
m841 470 466 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=3.609e-11 ps=1.77e-05 pd=3.577e-05 
+ nrs=0.05 nrd=0.14 
m842 469 287 470 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.008e-11 ad=1.36e-11 ps=3.81e-05 pd=1.77e-05 
+ nrs=0.12 nrd=0.05 
m843 471 290 469 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=3.5e-11 ps=4.183e-05 pd=6.21e-05 
+ nrs=0.06 nrd=0.04 
m844 1 466 471 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.938e-11 ad=4.62e-11 ps=6.998e-05 pd=4.183e-05 
+ nrs=0.08 nrd=0.06 
m845 471 287 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.938e-11 ps=4.183e-05 pd=6.998e-05 
+ nrs=0.06 nrd=0.08 
m846 0 469 468 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.609e-11 ad=3.008e-11 ps=3.577e-05 pd=3.81e-05 
+ nrs=0.14 nrd=0.12 
m847 472 397 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=3.609e-11 ps=1.77e-05 pd=3.577e-05 
+ nrs=0.05 nrd=0.14 
m848 468 290 472 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.008e-11 ad=1.36e-11 ps=3.81e-05 pd=1.77e-05 
+ nrs=0.12 nrd=0.05 
m849 473 469 468 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=3.5e-11 ps=4.183e-05 pd=6.21e-05 
+ nrs=0.06 nrd=0.04 
m850 1 397 473 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.938e-11 ad=4.62e-11 ps=6.998e-05 pd=4.183e-05 
+ nrs=0.08 nrd=0.06 
m851 473 290 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.938e-11 ps=4.183e-05 pd=6.998e-05 
+ nrs=0.06 nrd=0.08 
m852 474 476 475 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m853 0 392 474 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.609e-11 ad=2.507e-11 ps=3.577e-05 pd=2.557e-05 
+ nrs=0.14 nrd=0.1 
m854 474 369 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.609e-11 ps=2.557e-05 pd=3.577e-05 
+ nrs=0.1 nrd=0.14 
m855 475 476 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.938e-11 ps=3.13e-05 pd=6.998e-05 
+ nrs=0.06 nrd=0.08 
m856 477 392 475 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m857 1 369 477 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.938e-11 ad=4.62e-11 ps=6.998e-05 pd=3.13e-05 
+ nrs=0.08 nrd=0.06 
m858 0 390 478 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.895e-11 ad=2.562e-11 ps=1.878e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m859 1 390 478 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.308e-11 ad=2.694e-11 ps=3.899e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m860 0 480 479 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.895e-11 ad=2.562e-11 ps=1.878e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m861 1 480 479 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.308e-11 ad=2.694e-11 ps=3.899e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m862 0 403 481 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.895e-11 ad=2.562e-11 ps=1.878e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m863 1 403 481 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.308e-11 ad=2.694e-11 ps=3.899e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m864 482 478 464 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m865 0 332 482 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.609e-11 ad=1.36e-11 ps=3.577e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m866 464 478 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.969e-11 ps=1.73e-05 pd=3.499e-05 
+ nrs=0.12 nrd=0.15 
m867 1 332 464 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.969e-11 ad=2.31e-11 ps=3.499e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m868 483 392 476 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m869 0 369 483 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.609e-11 ad=1.36e-11 ps=3.577e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m870 476 392 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.969e-11 ps=1.73e-05 pd=3.499e-05 
+ nrs=0.12 nrd=0.15 
m871 1 369 476 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.969e-11 ad=2.31e-11 ps=3.499e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m872 484 481 480 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m873 0 326 484 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.609e-11 ad=1.36e-11 ps=3.577e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m874 480 481 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.969e-11 ps=1.73e-05 pd=3.499e-05 
+ nrs=0.12 nrd=0.15 
m875 1 326 480 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.969e-11 ad=2.31e-11 ps=3.499e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m876 485 487 486 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m877 0 479 485 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.609e-11 ad=2.507e-11 ps=3.577e-05 pd=2.557e-05 
+ nrs=0.14 nrd=0.1 
m878 485 488 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.609e-11 ps=2.557e-05 pd=3.577e-05 
+ nrs=0.1 nrd=0.14 
m879 486 487 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.938e-11 ps=3.13e-05 pd=6.998e-05 
+ nrs=0.06 nrd=0.08 
m880 489 479 486 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m881 1 488 489 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.938e-11 ad=4.62e-11 ps=6.998e-05 pd=3.13e-05 
+ nrs=0.08 nrd=0.06 
m882 0 306 488 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.895e-11 ad=2.562e-11 ps=1.878e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m883 1 306 488 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.308e-11 ad=2.694e-11 ps=3.899e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m884 0 424 487 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.895e-11 ad=2.562e-11 ps=1.878e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m885 1 424 487 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.308e-11 ad=2.694e-11 ps=3.899e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m886 0 486 490 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.895e-11 ad=2.562e-11 ps=1.878e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m887 1 486 490 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.308e-11 ad=2.694e-11 ps=3.899e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m888 491 493 492 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m889 0 311 491 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.609e-11 ad=2.507e-11 ps=3.577e-05 pd=2.557e-05 
+ nrs=0.14 nrd=0.1 
m890 491 238 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.609e-11 ps=2.557e-05 pd=3.577e-05 
+ nrs=0.1 nrd=0.14 
m891 492 493 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.938e-11 ps=3.13e-05 pd=6.998e-05 
+ nrs=0.06 nrd=0.08 
m892 494 311 492 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m893 1 238 494 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.938e-11 ad=4.62e-11 ps=6.998e-05 pd=3.13e-05 
+ nrs=0.08 nrd=0.06 
m894 495 311 493 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m895 0 238 495 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.609e-11 ad=1.36e-11 ps=3.577e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m896 493 311 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.969e-11 ps=1.73e-05 pd=3.499e-05 
+ nrs=0.12 nrd=0.15 
m897 1 238 493 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.969e-11 ad=2.31e-11 ps=3.499e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m898 496 498 497 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m899 0 316 496 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.609e-11 ad=2.507e-11 ps=3.577e-05 pd=2.557e-05 
+ nrs=0.14 nrd=0.1 
m900 496 490 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.609e-11 ps=2.557e-05 pd=3.577e-05 
+ nrs=0.1 nrd=0.14 
m901 497 498 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.938e-11 ps=3.13e-05 pd=6.998e-05 
+ nrs=0.06 nrd=0.08 
m902 499 316 497 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m903 1 490 499 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.938e-11 ad=4.62e-11 ps=6.998e-05 pd=3.13e-05 
+ nrs=0.08 nrd=0.06 
m904 500 70 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.804e-11 ps=1.13e-05 pd=1.788e-05 
+ nrs=0.21 nrd=0.28 
m905 0 490 500 0 nenh l=1.1e-06 w=8e-06 
+ as=1.804e-11 ad=1.32e-11 ps=1.788e-05 pd=1.13e-05 
+ nrs=0.28 nrd=0.21 
m906 501 70 500 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m907 1 490 501 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.938e-11 ad=2.38e-11 ps=6.998e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m908 502 503 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.804e-11 ps=1.13e-05 pd=1.788e-05 
+ nrs=0.21 nrd=0.28 
m909 0 70 502 0 nenh l=1.1e-06 w=8e-06 
+ as=1.804e-11 ad=1.32e-11 ps=1.788e-05 pd=1.13e-05 
+ nrs=0.28 nrd=0.21 
m910 504 503 502 1 penh l=1.1e-06 w=2.8e-05 
+ as=2.38e-11 ad=4.06e-11 ps=2.97e-05 pd=6.61e-05 
+ nrs=0.03 nrd=0.05 
m911 1 70 504 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.938e-11 ad=2.38e-11 ps=6.998e-05 pd=2.97e-05 
+ nrs=0.08 nrd=0.03 
m912 0 505 503 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.895e-11 ad=2.562e-11 ps=1.878e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m913 1 505 503 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.308e-11 ad=2.694e-11 ps=3.899e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m914 0 500 506 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.895e-11 ad=2.562e-11 ps=1.878e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m915 1 500 506 1 penh l=1.1e-06 w=1.56e-05 
+ as=3.308e-11 ad=2.694e-11 ps=3.899e-05 pd=3.57e-05 
+ nrs=0.14 nrd=0.11 
m916 507 316 498 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m917 0 490 507 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.609e-11 ad=1.36e-11 ps=3.577e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m918 498 316 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.969e-11 ps=1.73e-05 pd=3.499e-05 
+ nrs=0.12 nrd=0.15 
m919 1 490 498 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.969e-11 ad=2.31e-11 ps=3.499e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m920 508 83 505 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m921 0 490 508 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.609e-11 ad=1.36e-11 ps=3.577e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m922 505 83 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.969e-11 ps=1.73e-05 pd=3.499e-05 
+ nrs=0.12 nrd=0.15 
m923 1 490 505 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.969e-11 ad=2.31e-11 ps=3.499e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m924 509 506 510 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m925 0 83 509 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.609e-11 ad=1.36e-11 ps=3.577e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m926 510 506 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.969e-11 ps=1.73e-05 pd=3.499e-05 
+ nrs=0.12 nrd=0.15 
m927 1 83 510 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.969e-11 ad=2.31e-11 ps=3.499e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m928 0 415 411 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.609e-11 ad=3.008e-11 ps=3.577e-05 pd=3.81e-05 
+ nrs=0.14 nrd=0.12 
m929 511 510 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=3.609e-11 ps=1.77e-05 pd=3.577e-05 
+ nrs=0.05 nrd=0.14 
m930 411 413 511 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.008e-11 ad=1.36e-11 ps=3.81e-05 pd=1.77e-05 
+ nrs=0.12 nrd=0.05 
m931 512 415 411 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=3.5e-11 ps=4.183e-05 pd=6.21e-05 
+ nrs=0.06 nrd=0.04 
m932 1 510 512 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.938e-11 ad=4.62e-11 ps=6.998e-05 pd=4.183e-05 
+ nrs=0.08 nrd=0.06 
m933 512 413 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.938e-11 ps=4.183e-05 pd=6.998e-05 
+ nrs=0.06 nrd=0.08 
m934 513 413 339 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m935 0 502 513 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.609e-11 ad=2.507e-11 ps=3.577e-05 pd=2.557e-05 
+ nrs=0.14 nrd=0.1 
m936 513 415 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.609e-11 ps=2.557e-05 pd=3.577e-05 
+ nrs=0.1 nrd=0.14 
m937 339 413 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.938e-11 ps=3.13e-05 pd=6.998e-05 
+ nrs=0.06 nrd=0.08 
m938 514 502 339 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m939 1 415 514 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.938e-11 ad=4.62e-11 ps=6.998e-05 pd=3.13e-05 
+ nrs=0.08 nrd=0.06 
m940 515 416 516 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m941 0 413 515 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.609e-11 ad=1.36e-11 ps=3.577e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m942 516 416 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.969e-11 ps=1.73e-05 pd=3.499e-05 
+ nrs=0.12 nrd=0.15 
m943 1 413 516 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.969e-11 ad=2.31e-11 ps=3.499e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m944 517 519 518 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=2.8e-11 ps=2.557e-05 pd=3.81e-05 
+ nrs=0.1 nrd=0.11 
m945 0 502 517 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.609e-11 ad=2.507e-11 ps=3.577e-05 pd=2.557e-05 
+ nrs=0.14 nrd=0.1 
m946 517 516 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=2.507e-11 ad=3.609e-11 ps=2.557e-05 pd=3.577e-05 
+ nrs=0.1 nrd=0.14 
m947 518 519 1 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=5.938e-11 ps=3.13e-05 pd=6.998e-05 
+ nrs=0.06 nrd=0.08 
m948 520 502 518 1 penh l=1.1e-06 w=2.8e-05 
+ as=4.62e-11 ad=4.62e-11 ps=3.13e-05 pd=3.13e-05 
+ nrs=0.06 nrd=0.06 
m949 1 516 520 1 penh l=1.1e-06 w=2.8e-05 
+ as=5.938e-11 ad=4.62e-11 ps=6.998e-05 pd=3.13e-05 
+ nrs=0.08 nrd=0.06 
m950 521 510 519 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m951 0 516 521 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.609e-11 ad=1.36e-11 ps=3.577e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m952 519 510 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.969e-11 ps=1.73e-05 pd=3.499e-05 
+ nrs=0.12 nrd=0.15 
m953 1 516 519 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.969e-11 ad=2.31e-11 ps=3.499e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
m954 522 98 358 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.36e-11 ad=2.24e-11 ps=1.77e-05 pd=3.81e-05 
+ nrs=0.05 nrd=0.09 
m955 0 100 522 0 nenh l=1.1e-06 w=1.6e-05 
+ as=3.609e-11 ad=1.36e-11 ps=3.577e-05 pd=1.77e-05 
+ nrs=0.14 nrd=0.05 
m956 358 98 1 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.31e-11 ad=2.969e-11 ps=1.73e-05 pd=3.499e-05 
+ nrs=0.12 nrd=0.15 
m957 1 100 358 1 penh l=1.1e-06 w=1.4e-05 
+ as=2.969e-11 ad=2.31e-11 ps=3.499e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.12 
c0 285 0 9.3548e-14
c1 269 0 1.25582e-13
c2 206 0 9.0679e-14
c3 201 0 7.5745e-14
c4 151 0 1.72348e-13
c5 219 0 1.26195e-13
c6 449 0 1.4236e-14
c7 458 0 1.4236e-14
c8 432 0 1.1639e-13
c9 342 0 1.37304e-13
c10 437 0 1.17973e-13
c11 96 0 1.85078e-13
c12 420 0 1.30554e-13
c13 357 0 1.35189e-13
c14 256 0 1.38063e-13
c15 467 0 1.405e-14
c16 475 0 1.4236e-14
c17 492 0 1.4277e-14
c18 497 0 1.4236e-14
c19 518 0 1.4339e-14
c20 100 0 1.17274e-13
c21 98 0 1.07951e-13
c22 358 0 5.0945e-14
c23 1 0 3.69829e-13
c24 0 0 3.36103e-13
c29 516 0 4.7718e-14
c30 510 0 5.8123e-14
c31 519 0 3.0996e-14
c32 502 0 6.6827e-14
c33 517 0 9.87e-16
c34 413 0 7.3583e-14
c35 416 0 5.8642e-14
c36 415 0 5.4385e-14
c37 339 0 5.9788e-14
c38 513 0 9.87e-16
c39 512 0 1.101e-15
c40 411 0 5.5759e-14
c41 83 0 1.48914e-13
c42 506 0 2.8018e-14
c43 490 0 8.1293e-14
c44 505 0 4.562e-14
c45 316 0 6.2771e-14
c46 498 0 3.3153e-14
c47 500 0 4.5397e-14
c48 503 0 3.3078e-14
c49 70 0 1.24259e-13
c50 496 0 9.87e-16
c51 311 0 7.3166e-14
c52 493 0 3.8595e-14
c53 491 0 9.87e-16
c54 486 0 4.8188e-14
c55 424 0 4.1815e-14
c56 487 0 4.5024e-14
c57 306 0 4.8123e-14
c58 488 0 3.6561e-14
c59 479 0 3.5148e-14
c60 485 0 9.87e-16
c61 326 0 1.2196e-13
c62 480 0 3.8046e-14
c63 369 0 1.50624e-13
c64 392 0 5.7751e-14
c65 476 0 4.1331e-14
c66 464 0 7.1094e-14
c67 403 0 3.6552e-14
c68 481 0 3.4107e-14
c69 390 0 3.6511e-14
c70 478 0 3.8907e-14
c71 474 0 9.87e-16
c72 290 0 6.424e-14
c73 473 0 1.101e-15
c74 397 0 2.51985e-13
c75 469 0 3.6589e-14
c76 287 0 9.0004e-14
c77 471 0 1.101e-15
c78 466 0 2.8688e-14
c79 468 0 3.8204e-14
c80 381 0 7.0837e-14
c81 384 0 6.9789e-14
c82 459 0 4.3045e-14
c83 454 0 2.4007e-14
c84 447 0 5.848e-14
c85 450 0 4.333e-14
c86 461 0 9.87e-16
c87 386 0 7.7514e-14
c88 457 0 9.87e-16
c89 363 0 7.8445e-14
c90 455 0 3.2446e-14
c91 373 0 5.796e-14
c92 364 0 8.6993e-14
c93 445 0 5.1892e-14
c94 275 0 7.393e-14
c95 452 0 9.87e-16
c96 395 0 6.3633e-14
c97 448 0 9.87e-16
c98 443 0 2.5922e-14
c99 441 0 9.917e-14
c100 440 0 9.9771e-14
c101 281 0 5.5115e-14
c102 362 0 4.0274e-14
c103 267 0 5.8232e-14
c104 372 0 4.2339e-14
c105 380 0 3.737e-14
c106 389 0 3.8526e-14
c107 394 0 4.5735e-14
c108 247 0 8.1498e-14
c109 427 0 4.8452e-14
c110 409 0 4.6692e-14
c111 414 0 4.3822e-14
c112 192 0 7.4841e-14
c113 288 0 1.0289e-13
c114 348 0 5.3424e-14
c115 406 0 3.9672e-14
c116 387 0 3.6204e-14
c117 304 0 7.5166e-14
c118 417 0 1.80597e-13
c119 429 0 3.532e-14
c120 407 0 3.527e-14
c121 435 0 3.9626e-14
c122 366 0 2.9532e-14
c123 370 0 3.1301e-14
c124 371 0 2.5521e-14
c125 404 0 2.6087e-14
c126 408 0 2.4172e-14
c127 418 0 1.74391e-13
c128 436 0 9.87e-16
c129 250 0 4.8292e-14
c130 431 0 9.87e-16
c131 313 0 3.4301e-14
c132 428 0 9.87e-16
c133 423 0 9.87e-16
c134 324 0 9.9186e-14
c135 1 0 4.09593e-13
c136 0 0 3.56977e-13
c138 260 0 5.4138e-14
c139 318 0 7.404e-14
c140 347 0 3.6135e-14
c141 336 0 4.9514e-14
c142 225 0 7.7131e-14
c143 405 0 3.1013e-14
c144 385 0 2.3946e-14
c145 399 0 9.87e-16
c146 293 0 8.2559e-14
c147 398 0 1.101e-15
c148 57 0 8.2694e-14
c149 298 0 1.19246e-13
c150 378 0 9.026e-14
c151 332 0 8.4573e-14
c152 377 0 4.7252e-14
c153 330 0 7.3016e-14
c154 368 0 1.101e-15
c155 274 0 6.6559e-14
c156 271 0 5.6973e-14
c157 265 0 3.8128e-14
c158 279 0 4.9192e-14
c159 282 0 1.0465e-13
c160 295 0 9.9094e-14
c161 291 0 3.2976e-14
c162 283 0 1.08879e-13
c163 294 0 1.3075e-13
c164 297 0 3.192e-14
c165 300 0 1.2631e-13
c166 303 0 4.2247e-14
c167 299 0 1.19665e-13
c168 307 0 5.2382e-14
c169 315 0 2.9448e-14
c170 320 0 1.30165e-13
c171 337 0 2.8393e-14
c172 319 0 1.9552e-13
c173 309 0 5.6436e-14
c174 343 0 3.1087e-14
c175 353 0 1.10098e-13
c176 351 0 3.2125e-14
c177 173 0 1.54035e-13
c178 286 0 5.9742e-14
c179 352 0 1.30832e-13
c180 344 0 6.1676e-14
c181 273 0 3.1472e-14
c182 277 0 3.0126e-14
c183 302 0 2.5542e-14
c184 361 0 1.101e-15
c185 181 0 5.071e-14
c186 234 0 8.9161e-14
c187 261 0 3.2903e-14
c188 1 0 3.89672e-13
c189 186 0 4.8195e-14
c190 0 0 3.47231e-13
c191 86 0 7.3653e-14
c192 356 0 9.87e-16
c193 350 0 9.87e-16
c194 346 0 9.87e-16
c195 341 0 9.87e-16
c196 340 0 1.101e-15
c197 231 0 5.3145e-14
c198 270 0 2.6827e-14
c199 310 0 3.4815e-14
c200 175 0 9.4739e-14
c201 249 0 3.819e-14
c202 124 0 4.8585e-14
c203 223 0 9.2037e-14
c204 113 0 1.04194e-13
c205 268 0 9.87e-16
c206 3 0 9.6985e-14
c207 101 0 5.1031e-14
c208 12 0 7.2011e-14
c209 264 0 9.87e-16
c210 229 0 3.1119e-14
c211 149 0 8.0471e-14
c212 242 0 4.6516e-14
c213 185 0 6.0641e-14
c214 257 0 3.109e-14
c215 188 0 4.1948e-14
c216 198 0 3.7663e-14
c217 193 0 1.13373e-13
c218 230 0 4.6003e-14
c219 182 0 6.7499e-14
c220 179 0 6.3804e-14
c221 235 0 3.4856e-14
c222 189 0 2.7822e-14
c223 237 0 3.1267e-14
c224 240 0 3.2488e-14
c225 241 0 2.4869e-14
c226 263 0 1.101e-15
c227 184 0 8.4766e-14
c228 1 0 4.20533e-13
c229 0 0 3.66328e-13
c231 255 0 9.87e-16
c232 252 0 1.101e-15
c233 143 0 8.96e-14
c234 139 0 3.4758e-14
c235 140 0 5.5405e-14
c236 109 0 2.067e-13
c237 169 0 2.7477e-14
c238 162 0 1.0615e-13
c239 238 0 1.26271e-13
c240 157 0 6.4542e-14
c241 227 0 8.8673e-14
c242 226 0 8.9349e-14
c243 155 0 5.2587e-14
c244 214 0 6.5121e-14
c245 221 0 3.0702e-14
c246 19 0 1.16853e-13
c247 137 0 4.6969e-14
c248 135 0 4.8261e-14
c249 217 0 3.7383e-14
c250 218 0 9.87e-16
c251 132 0 4.9809e-14
c252 50 0 7.938e-14
c253 212 0 2.9068e-14
c254 210 0 3.1001e-14
c255 203 0 1.1088e-13
c256 115 0 5.719e-14
c257 207 0 4.0153e-14
c258 205 0 9.87e-16
c259 48 0 9.7985e-14
c260 195 0 4.6287e-14
c261 119 0 3.6725e-14
c262 197 0 3.1282e-14
c263 200 0 9.87e-16
c264 196 0 9.87e-16
c265 105 0 3.0823e-14
c266 107 0 7.041e-14
c267 111 0 7.5815e-14
c268 114 0 1.728e-13
c269 121 0 8.9374e-14
c270 145 0 9.4937e-14
c271 144 0 1.1127e-13
c272 106 0 2.4869e-14
c273 161 0 9.2391e-14
c274 183 0 9.87e-16
c275 1 0 4.19137e-13
c276 0 0 3.65972e-13
c279 171 0 2.6055e-14
c280 164 0 1.18876e-13
c281 163 0 5.1009e-14
c282 159 0 5.3353e-14
c283 158 0 9.959e-14
c284 166 0 3.8136e-14
c285 170 0 4.4244e-14
c286 167 0 2.22661e-13
c287 65 0 4.5224e-14
c288 81 0 3.7402e-14
c289 64 0 2.8731e-14
c290 75 0 5.3295e-14
c291 152 0 3.086e-14
c292 154 0 9.87e-16
c293 76 0 3.8882e-14
c294 150 0 9.87e-16
c295 35 0 6.0375e-14
c296 142 0 4.2156e-14
c297 62 0 4.6971e-14
c298 133 0 2.8045e-14
c299 34 0 6.8054e-14
c300 136 0 9.87e-16
c301 28 0 9.1259e-14
c302 129 0 3.8544e-14
c303 130 0 1.101e-15
c304 125 0 3.1613e-14
c305 127 0 1.101e-15
c306 110 0 6.771e-14
c307 14 0 7.0937e-14
c308 122 0 1.101e-15
c309 7 0 1.07025e-13
c310 24 0 8.8434e-14
c311 104 0 4.986e-14
c312 116 0 7.208e-14
c313 102 0 3.3138e-14
c314 44 0 5.7068e-14
c315 25 0 6.7516e-14
c316 23 0 3.2865e-14
c317 46 0 1.10673e-13
c318 36 0 3.1073e-14
c319 30 0 6.9429e-14
c320 58 0 5.8471e-14
c321 8 0 3.3422e-14
c322 27 0 4.2663e-14
c323 17 0 3.7922e-14
c324 37 0 3.5949e-14
c325 60 0 2.5963e-14
c326 85 0 1.26819e-13
c327 53 0 1.55534e-13
c328 94 0 3.4604e-14
c329 1 0 4.20805e-13
c330 0 0 3.6679e-13
c334 87 0 4.8219e-14
c335 89 0 4.3705e-14
c336 95 0 1.101e-15
c337 68 0 5.8667e-14
c338 90 0 3.4997e-14
c339 92 0 1.101e-15
c340 78 0 7.595e-14
c341 84 0 9.87e-16
c342 72 0 3.2614e-14
c343 71 0 3.109e-14
c344 61 0 4.5029e-14
c345 79 0 1.101e-15
c346 39 0 1.08107e-13
c347 67 0 2.6786e-14
c348 55 0 1.02787e-13
c349 15 0 1.54841e-13
c350 56 0 9.87e-16
c351 41 0 3.0966e-14
c352 40 0 3.1526e-14
c353 21 0 3.5197e-14
c354 20 0 3.7032e-14
c355 32 0 3.4338e-14
c356 31 0 3.1586e-14
c357 16 0 2.8851e-14
c358 9 0 3.4364e-14
c359 5 0 4.304e-14
c360 4 0 4.0186e-14
c361 170 114 9.74e-16
c362 311 407 1.58e-16
c363 110 4 1.58e-16
c364 432 326 1.58e-16
c365 173 233 1.926e-15
c366 510 1 8.959e-15
c367 516 0 5.333e-15
c368 119 107 1.58e-16
c369 50 109 1.58e-16
c370 1 313 1.862e-15
c371 397 332 3.15e-16
c372 48 30 1.58e-16
c373 83 161 1.58e-16
c374 353 1 8.3e-16
c375 1 404 3.815e-15
c376 76 114 1.58e-16
c377 225 1 6.989e-15
c378 502 503 8.89e-16
c379 1 142 5.854e-15
c380 28 30 1.58e-16
c381 227 46 1.58e-16
c382 0 27 3.719e-15
c383 100 184 1.58e-16
c384 256 0 1.327e-15
c385 285 1 8.3e-16
c386 300 223 1.58e-16
c387 254 0 8.06e-16
c388 350 0 2.893e-15
c389 386 288 3.15e-16
c390 447 364 1.58e-16
c391 450 373 3.15e-16
c392 151 293 3.15e-16
c393 420 510 4.73e-16
c394 336 319 1.132e-15
c395 0 461 2.893e-15
c396 326 332 3.15e-16
c397 80 0 8.06e-16
c398 361 173 9.54e-16
c399 86 78 2.02e-16
c400 353 55 1.58e-16
c401 432 311 1.58e-16
c402 68 53 4.73e-16
c403 176 0 8.06e-16
c404 1 299 3.724e-15
c405 369 478 3.15e-16
c406 392 390 2.22e-16
c407 479 397 3.15e-16
c408 164 35 3.15e-16
c409 227 1 8.3e-16
c410 86 0 8.3e-16
c411 282 110 4.73e-16
c412 344 343 2.848e-15
c413 227 144 1.58e-16
c414 353 75 1.58e-16
c415 218 0 2.893e-15
c416 96 464 1.58e-16
c417 192 274 3.54e-16
c418 397 472 4.8e-16
c419 100 356 6.62e-16
c420 300 107 1.58e-16
c421 299 114 1.58e-16
c422 57 227 1.58e-16
c423 96 214 1.58e-16
c424 304 238 1.58e-16
c425 1 145 4.761e-15
c426 299 207 1.58e-16
c427 96 352 1.58e-16
c428 301 299 1.926e-15
c429 326 479 1.58e-16
c430 19 227 3.15e-16
c431 33 1 8.06e-16
c432 81 1 1.301e-15
c433 193 119 1.58e-16
c434 125 1 3.189e-15
c435 295 1 8.3e-16
c436 50 7 1.58e-16
c437 250 1 1.327e-15
c438 109 143 1.58e-16
c439 320 0 8.3e-16
c440 70 0 1.612e-15
c441 0 508 8.06e-16
c442 15 35 3.15e-16
c443 0 183 2.893e-15
c444 304 249 7.32e-16
c445 0 500 3.719e-15
c446 424 1 3.293e-15
c447 62 0 1.612e-15
c448 330 286 1.58e-16
c449 466 287 1.58e-16
c450 0 203 1.0423e-14
c451 274 273 7.32e-16
c452 0 367 8.06e-16
c453 419 417 1.926e-15
c454 169 1 1.862e-15
c455 70 503 1.323e-15
c456 151 288 3.15e-16
c457 357 247 1.58e-16
c458 253 0 8.06e-16
c459 258 1 1.565e-15
c460 50 0 1.327e-15
c461 96 1 8.3e-16
c462 324 298 6.3e-16
c463 70 418 1.58e-16
c464 0 407 3.194e-15
c465 269 0 8.3e-16
c466 206 1 8.3e-16
c467 353 167 1.58e-16
c468 162 319 1.58e-16
c469 1 373 1.327e-15
c470 77 0 8.06e-16
c471 0 277 2.877e-15
c472 164 15 1.58e-16
c473 37 46 3.15e-16
c474 417 132 2.06e-16
c475 1 441 4.761e-15
c476 0 446 8.06e-16
c477 96 114 1.58e-16
c478 256 225 5.74e-16
c479 418 158 1.58e-16
c480 519 516 1.58e-16
c481 416 1 1.862e-15
c482 413 0 5.868e-15
c483 402 0 8.06e-16
c484 226 114 1.58e-16
c485 219 167 6.3e-16
c486 70 0 8.3e-16
c487 513 415 6.62e-16
c488 295 1 8.3e-16
c489 332 0 1.327e-15
c490 348 346 6.62e-16
c491 17 16 1.723e-15
c492 231 0 3.724e-15
c493 330 279 4.73e-16
c494 397 394 4.73e-16
c495 287 386 3.15e-16
c496 227 167 1.58e-16
c497 1 37 4.761e-15
c498 256 1 8.3e-16
c499 432 0 1.327e-15
c500 279 223 7.32e-16
c501 50 20 9.74e-16
c502 381 1 5.841e-15
c503 306 486 1.9e-16
c504 0 390 1.827e-15
c505 1 478 3.163e-15
c506 141 39 1.926e-15
c507 169 1 1.301e-15
c508 143 149 6.3e-16
c509 65 164 1.58e-16
c510 238 1 2.247e-15
c511 423 304 6.36e-16
c512 339 348 1.58e-16
c513 363 288 3.15e-16
c514 447 448 6.62e-16
c515 420 416 1.58e-16
c516 418 332 3.15e-16
c517 505 397 3.15e-16
c518 22 20 1.926e-15
c519 109 144 3.15e-16
c520 66 1 8.06e-16
c521 1 232 8.06e-16
c522 341 343 1.042e-15
c523 18 16 1.926e-15
c524 113 203 1.58e-16
c525 93 0 8.06e-16
c526 392 397 4.73e-16
c527 26 1 8.06e-16
c528 57 109 1.58e-16
c529 1 339 3.293e-15
c530 21 0 3.756e-15
c531 35 53 3.15e-16
c532 319 283 1.58e-16
c533 83 319 1.58e-16
c534 256 175 3.15e-16
c535 420 478 3.15e-16
c536 357 390 1.58e-16
c537 508 83 7.96e-16
c538 83 500 3.15e-16
c539 0 487 2.912e-15
c540 251 0 8.06e-16
c541 0 332 3.689e-15
c542 12 105 4.6e-16
c543 169 234 1.58e-16
c544 249 1 1.862e-15
c545 109 19 1.58e-16
c546 304 427 1.58e-16
c547 195 196 1.042e-15
c548 300 17 3.15e-16
c549 24 110 3.15e-16
c550 420 339 1.58e-16
c551 164 34 3.34e-16
c552 283 3 3.15e-16
c553 186 0 8.3e-16
c554 299 116 1.58e-16
c555 151 212 1.58e-16
c556 275 0 3.474e-15
c557 30 25 1.58e-16
c558 164 53 3.15e-16
c559 294 197 3.15e-16
c560 83 159 1.74e-16
c561 188 195 1.58e-16
c562 437 306 1.58e-16
c563 7 46 3.15e-16
c564 353 0 8.3e-16
c565 294 15 1.58e-16
c566 290 378 1.58e-16
c567 193 5 1.58e-16
c568 418 1 8.3e-16
c569 203 48 1.275e-15
c570 20 21 1.88e-15
c571 298 281 1.58e-16
c572 70 85 1.58e-16
c573 151 287 3.15e-16
c574 432 406 3.15e-16
c575 14 0 3.689e-15
c576 28 25 3.15e-16
c577 149 144 9.74e-16
c578 0 209 8.06e-16
c579 0 46 5.051e-15
c580 1 36 3.724e-15
c581 219 0 1.327e-15
c582 299 223 1.58e-16
c583 256 86 1.58e-16
c584 1 119 1.862e-15
c585 0 195 5.051e-15
c586 7 1 5.437e-15
c587 467 0 1.05e-15
c588 475 1 3.293e-15
c589 158 85 3.39e-16
c590 63 61 1.926e-15
c591 7 144 1.58e-16
c592 0 275 8.3e-16
c593 0 459 3.189e-15
c594 0 227 3.756e-15
c595 61 0 2.771e-15
c596 353 155 1.58e-16
c597 15 34 1.58e-16
c598 385 1 5.001e-15
c599 484 481 7.96e-16
c600 320 235 3.15e-16
c601 15 53 1.58e-16
c602 63 1 8.06e-16
c603 186 0 1.862e-15
c604 520 502 3.306e-15
c605 109 167 1.578e-15
c606 348 417 1.58e-16
c607 144 0 8.3e-16
c608 353 0 8.3e-16
c609 175 253 7.96e-16
c610 411 438 3.306e-15
c611 299 107 1.58e-16
c612 418 1 8.3e-16
c613 1 278 8.06e-16
c614 7 19 3.15e-16
c615 269 386 3.15e-16
c616 1 121 1.2359e-14
c617 57 0 1.327e-15
c618 14 111 3.15e-16
c619 328 294 7.96e-16
c620 329 297 7.96e-16
c621 14 30 4.6e-16
c622 151 157 3.15e-16
c623 212 50 6.54e-16
c624 0 397 1.862e-15
c625 1 469 3.189e-15
c626 485 487 1.042e-15
c627 217 1 4.591e-15
c628 155 227 3.15e-16
c629 55 0 7.16e-15
c630 0 234 2.683e-15
c631 119 1 1.327e-15
c632 65 53 7.32e-16
c633 19 0 3.719e-15
c634 150 152 1.042e-15
c635 300 1 8.3e-16
c636 316 427 1.58e-16
c637 1 309 5.677e-15
c638 476 332 1.58e-16
c639 227 0 8.3e-16
c640 129 1 7.098e-15
c641 75 0 1.327e-15
c642 96 223 1.58e-16
c643 502 415 4.82e-16
c644 20 1 3.724e-15
c645 237 242 1.46e-16
c646 478 464 1.132e-15
c647 420 469 1.58e-16
c648 357 397 3.15e-16
c649 319 230 3.15e-16
c650 505 503 1.58e-16
c651 0 326 2.144e-15
c652 332 286 3.15e-16
c653 428 313 6.36e-16
c654 113 227 1.58e-16
c655 206 1 8.3e-16
c656 1 101 1.862e-15
c657 149 167 1.58e-16
c658 260 1 1.327e-15
c659 352 39 1.58e-16
c660 151 319 1.58e-16
c661 1 414 4.616e-15
c662 0 394 5.338e-15
c663 452 445 1.042e-15
c664 98 185 1.58e-16
c665 250 162 1.58e-16
c666 441 1 8.3e-16
c667 357 250 1.58e-16
c668 83 81 1.58e-16
c669 19 20 7.32e-16
c670 357 326 1.58e-16
c671 521 0 8.06e-16
c672 294 4 1.58e-16
c673 282 15 1.58e-16
c674 206 207 2.69e-15
c675 300 1 8.3e-16
c676 219 285 1.58e-16
c677 201 206 4.73e-16
c678 0 382 8.06e-16
c679 151 269 3.15e-16
c680 206 12 3.15e-16
c681 0 311 4.462e-15
c682 392 0 1.892e-15
c683 469 290 6.69e-16
c684 227 30 1.58e-16
c685 143 235 1.263e-15
c686 338 0 8.06e-16
c687 101 44 7.32e-16
c688 195 48 3.15e-16
c689 109 0 2.441e-15
c690 100 1 8.3e-16
c691 206 440 1.58e-16
c692 201 441 1.58e-16
c693 336 0 3.189e-15
c694 219 1 8.3e-16
c695 441 12 1.58e-16
c696 347 1 1.327e-15
c697 1 403 3.289e-15
c698 76 158 1.58e-16
c699 450 445 1.58e-16
c700 447 275 1.58e-16
c701 441 44 1.58e-16
c702 175 353 1.58e-16
c703 83 397 3.15e-16
c704 163 1 3.724e-15
c705 400 386 3.306e-15
c706 440 441 2.068e-15
c707 1 460 1.565e-15
c708 79 1 3.083e-15
c709 1 233 8.06e-16
c710 247 320 1.58e-16
c711 336 418 1.58e-16
c712 339 409 6.17e-16
c713 357 311 1.58e-16
c714 89 0 4.303e-15
c715 1 307 6.289e-15
c716 227 28 1.58e-16
c717 324 0 1.327e-15
c718 339 1 4.533e-15
c719 133 0 2.912e-15
c720 181 185 1.58e-16
c721 114 39 1.58e-16
c722 1 85 1.301e-15
c723 418 137 1.58e-16
c724 306 247 1.58e-16
c725 326 281 1.58e-16
c726 137 121 2.02e-16
c727 282 294 1.58e-16
c728 319 320 2.049e-15
c729 304 417 1.58e-16
c730 369 455 1.58e-16
c731 420 403 1.58e-16
c732 0 106 2.493e-15
c733 110 114 9.74e-16
c734 126 121 4.8e-16
c735 132 34 4.6e-16
c736 83 250 3.15e-16
c737 324 418 7.31e-16
c738 109 155 1.58e-16
c739 1 276 8.06e-16
c740 347 349 3.306e-15
c741 387 389 1.58e-16
c742 269 363 3.15e-16
c743 336 0 1.827e-15
c744 55 79 9.54e-16
c745 12 110 1.58e-16
c746 461 454 6.62e-16
c747 342 344 1.58e-16
c748 62 58 1.58e-16
c749 319 104 1.58e-16
c750 519 397 3.15e-16
c751 109 0 5.163e-15
c752 249 229 1.132e-15
c753 110 44 1.58e-16
c754 100 1 8.3e-16
c755 260 234 6.73e-16
c756 339 318 1.58e-16
c757 255 185 6.36e-16
c758 269 270 2.69e-15
c759 440 110 1.58e-16
c760 275 279 6.17e-16
c761 0 324 3.724e-15
c762 0 149 5.833e-15
c763 0 439 8.06e-16
c764 493 238 1.58e-16
c765 109 113 1.59e-15
c766 104 3 1.58e-16
c767 437 435 3.005e-15
c768 469 464 3.15e-16
c769 0 503 2.493e-15
c770 417 214 1.58e-16
c771 139 1 2.514e-15
c772 342 288 3.15e-16
c773 397 386 3.6e-16
c774 143 157 1.686e-15
c775 332 299 9.74e-16
c776 417 352 3.15e-16
c777 98 181 1.58e-16
c778 100 234 1.58e-16
c779 162 0 3.439e-15
c780 357 0 1.327e-15
c781 449 0 1.327e-15
c782 458 1 3.293e-15
c783 217 137 1.96e-16
c784 256 353 1.614e-15
c785 441 364 3.15e-16
c786 193 105 1.58e-16
c787 96 70 5.48e-16
c788 302 303 1.46e-16
c789 357 418 1.58e-16
c790 392 476 1.36e-15
c791 186 183 6.62e-16
c792 155 149 1.147e-15
c793 109 111 1.58e-16
c794 1 442 8.06e-16
c795 502 510 3.15e-16
c796 515 0 8.06e-16
c797 96 432 1.58e-16
c798 149 0 1.327e-15
c799 109 48 3.15e-16
c800 96 158 1.58e-16
c801 417 1 8.3e-16
c802 170 1 5.854e-15
c803 357 0 8.3e-16
c804 167 161 3.15e-16
c805 81 80 7.96e-16
c806 109 28 5.27e-16
c807 24 15 4.73e-16
c808 306 487 1.74e-16
c809 7 0 4.295e-15
c810 139 1 1.301e-15
c811 281 0 1.892e-15
c812 316 417 1.58e-16
c813 411 435 3.54e-16
c814 73 1 8.06e-16
c815 234 361 3.137e-15
c816 1 455 3.189e-15
c817 299 1 8.3e-16
c818 417 114 1.58e-16
c819 1 425 1.565e-15
c820 76 1 1.862e-15
c821 78 0 5.051e-15
c822 83 0 1.827e-15
c823 0 283 3.756e-15
c824 140 223 9.74e-16
c825 1 512 3.083e-15
c826 369 389 1.58e-16
c827 175 109 1.58e-16
c828 318 417 3.15e-16
c829 1 374 8.06e-16
c830 45 16 7.96e-16
c831 83 418 1.58e-16
c832 269 267 4.73e-16
c833 432 238 1.58e-16
c834 67 69 1.926e-15
c835 12 194 7.96e-16
c836 320 145 1.58e-16
c837 62 145 1.58e-16
c838 116 110 5.55e-16
c839 363 459 1.58e-16
c840 184 263 6.36e-16
c841 151 295 1.58e-16
c842 269 271 2.02e-16
c843 1 372 5.854e-15
c844 0 281 3.439e-15
c845 440 362 1.58e-16
c846 445 373 1.96e-16
c847 210 1 4.616e-15
c848 124 294 1.58e-16
c849 58 46 1.96e-16
c850 0 241 2.493e-15
c851 1 453 1.565e-15
c852 7 111 3.15e-16
c853 151 326 2.06e-16
c854 7 30 3.15e-16
c856 83 0 8.3e-16
c857 0 434 8.06e-16
c858 299 1 8.3e-16
c859 319 1 8.3e-16
c860 410 348 1.926e-15
c861 185 187 3.306e-15
c862 61 58 7.32e-16
c863 57 247 1.58e-16
c864 342 287 3.15e-16
c865 162 163 7.32e-16
c866 7 48 1.58e-16
c867 289 287 1.926e-15
c868 314 1 8.06e-16
c869 227 25 1.58e-16
c870 111 0 8.3e-16
c871 1 58 6.478e-15
c872 0 30 2.912e-15
c873 96 1 8.3e-16
c874 159 61 1.58e-16
c875 7 28 1.263e-15
c876 109 86 3.15e-16
c877 57 319 1.58e-16
c878 0 476 3.189e-15
c879 226 1 3.724e-15
c880 285 293 3.15e-16
c881 98 1 1.862e-15
c882 100 0 2.144e-15
c883 3 1 1.327e-15
c884 159 1 8.3e-16
c885 48 0 1.327e-15
c886 352 164 1.58e-16
c887 0 447 5.051e-15
c888 1 236 8.06e-16
c889 57 58 2.02e-16
c890 198 196 6.36e-16
c891 293 1 1.862e-15
c892 306 397 3.47e-16
c893 64 85 1.58e-16
c894 28 0 2.771e-15
c896 231 249 3.15e-16
c897 321 1 8.06e-16
c898 344 337 2.6e-16
c899 352 351 1.171e-15
c900 416 502 1.58e-16
c901 324 279 1.58e-16
c902 357 476 3.15e-16
c903 250 320 1.58e-16
c904 308 307 1.926e-15
c905 100 357 1.58e-16
c906 98 420 1.58e-16
c907 19 115 1.58e-16
c908 198 188 1.03e-16
c909 274 1 3.724e-15
c910 363 365 1.926e-15
c911 159 55 3.15e-16
c912 75 58 1.58e-16
c913 35 114 3.15e-16
c914 157 167 1.58e-16
c915 454 459 4.39e-16
c916 1 105 2.514e-15
c917 238 1 4.761e-15
c918 373 372 1.58e-16
c919 489 479 3.306e-15
c920 96 1 8.3e-16
c921 206 193 3.15e-16
c922 192 1 8.3e-16
c923 386 0 4.492e-15
c924 155 156 3.306e-15
c925 0 235 2.493e-15
c926 79 78 6.36e-16
c927 83 163 3.15e-16
c928 226 1 8.3e-16
c929 143 145 1.58e-16
c930 90 68 1.275e-15
c931 352 15 1.58e-16
c932 0 198 4.492e-15
c933 71 0 3.306e-15
c934 212 0 2.912e-15
c935 441 193 3.15e-16
c936 0 343 3.189e-15
c937 1 351 4.591e-15
c938 70 427 1.58e-16
c939 83 85 1.58e-16
c940 296 294 1.926e-15
c941 502 339 2.02e-16
c942 0 161 7.199e-15
c943 164 114 3.15e-16
c944 175 310 1.58e-16
c945 507 316 7.96e-16
c946 1 369 8.461e-15
c947 0 484 8.06e-16
c948 249 1 2.565e-15
c949 201 192 1.58e-16
c950 342 247 1.58e-16
c951 192 12 1.58e-16
c952 151 0 8.3e-16
c953 311 306 1.58e-16
c954 319 167 1.58e-16
c955 413 435 3.15e-16
c957 440 192 1.58e-16
c958 1 288 3.724e-15
c959 24 282 1.58e-16
c960 145 46 1.58e-16
c961 1 273 4.616e-15
c962 105 1 1.301e-15
c963 294 214 1.58e-16
c964 1 15 2.247e-15
c965 417 330 1.58e-16
c966 151 418 1.58e-16
c967 52 36 7.96e-16
c968 86 0 2.6e-15
c969 420 369 3.15e-16
c970 417 223 1.58e-16
c971 109 203 1.58e-16
c972 283 5 1.58e-16
c973 269 167 1.58e-16
c974 267 375 7.96e-16
c975 369 384 3.15e-16
c976 397 429 3.15e-16
c977 256 468 1.58e-16
c978 264 12 1.042e-15
c979 15 114 1.58e-16
c980 201 197 2.69e-15
c981 145 1 8.3e-16
c982 207 15 1.58e-16
c983 151 0 8.3e-16
c984 437 1 3.293e-15
c985 81 61 9.74e-16
c986 144 145 2.049e-15
c987 52 0 8.06e-16
c988 424 486 3.34e-16
c989 380 281 1.58e-16
c990 250 143 3.54e-16
c991 231 309 4.48e-16
c992 81 1 1.862e-15
c993 57 145 1.58e-16
c994 444 440 7.96e-16
c995 76 64 1.58e-16
c996 0 157 1.612e-15
c997 341 337 6.36e-16
c998 440 442 1.926e-15
c999 352 53 1.58e-16
c1000 93 94 4.8e-16
c1001 1 294 3.724e-15
c1002 0 320 3.756e-15
c1003 369 290 1.58e-16
c1004 0 9 3.756e-15
c1005 342 298 3.15e-16
c1006 0 415 4.545e-15
c1007 270 0 3.189e-15
c1008 135 121 1.88e-16
c1009 65 114 1.58e-16
c1010 306 0 1.892e-15
c1011 432 478 3.15e-16
c1012 418 320 1.58e-16
c1013 433 250 3.306e-15
c1014 320 121 1.58e-16
c1015 151 217 3.15e-16
c1016 158 39 1.58e-16
c1017 295 46 1.58e-16
c1018 81 55 4.6e-16
c1019 137 226 1.58e-16
c1020 294 207 3.15e-16
c1021 306 418 1.58e-16
c1022 386 447 1.58e-16
c1023 457 459 1.042e-15
c1024 247 0 1.327e-15
c1025 151 300 1.58e-16
c1026 96 324 1.58e-16
c1027 480 326 1.58e-16
c1028 110 123 7.96e-16
c1029 127 125 3.137e-15
c1030 294 12 1.58e-16
c1031 363 0 2.771e-15
c1032 50 121 1.58e-16
c1033 155 157 3.15e-16
c1034 3 188 1.58e-16
c1035 165 1 8.06e-16
c1036 198 48 7.32e-16
c1037 294 44 1.58e-16
c1038 332 378 3.15e-16
c1039 437 424 1.58e-16
c1040 7 25 1.578e-15
c1041 319 0 8.3e-16
c1042 440 294 1.58e-16
c1043 0 522 8.06e-16
c1044 411 1 3.724e-15
c1045 320 129 1.58e-16
c1046 478 332 4.48e-16
c1047 157 0 3.719e-15
c1048 132 214 3.15e-16
c1049 295 1 8.3e-16
c1051 285 287 3.15e-16
c1052 306 0 8.3e-16
c1053 369 395 1.58e-16
c1054 34 114 1.58e-16
c1055 295 144 1.58e-16
c1056 0 115 4.462e-15
c1057 114 53 3.15e-16
c1058 0 25 5.331e-15
c1059 140 1 1.862e-15
c1060 98 171 9.74e-16
c1061 206 1 3.293e-15
c1062 101 1 3.289e-15
c1063 3 0 1.612e-15
c1064 143 232 1.926e-15
c1065 175 235 3.15e-16
c1066 287 1 5.151e-15
c1067 98 1 8.3e-16
c1068 381 288 1.58e-16
c1069 1 204 8.06e-16
c1070 231 307 9.74e-16
c1071 96 0 8.3e-16
c1072 420 1 8.3e-16
c1073 217 135 4.41e-16
c1074 456 363 1.926e-15
c1075 109 353 1.58e-16
c1076 441 1 8.3e-16
c1077 330 274 3.15e-16
c1078 326 57 3.66e-16
c1079 1 384 6.214e-15
c1080 167 145 3.15e-16
c1081 369 464 1.58e-16
c1082 86 161 1.58e-16
c1083 1 94 7.098e-15
c1084 182 185 1.58e-16
c1085 1 6 8.06e-16
c1086 173 185 3.15e-16
c1087 352 242 1.58e-16
c1088 319 0 8.3e-16
c1089 215 212 7.96e-16
c1090 397 435 3.15e-16
c1091 256 437 1.58e-16
c1092 275 378 3.15e-16
c1093 437 381 3.15e-16
c1094 342 459 1.58e-16
c1095 269 450 3.15e-16
c1096 333 0 8.06e-16
c1097 228 226 1.926e-15
c1098 151 286 1.58e-16
c1099 115 0 1.892e-15
c1100 319 113 1.58e-16
c1101 109 227 1.58e-16
c1102 96 64 1.58e-16
c1103 358 397 3.15e-16
c1104 1 290 3.724e-15
c1105 159 78 1.58e-16
c1106 12 4 9.74e-16
c1107 140 1 3.189e-15
c1108 267 0 1.05e-15
c1109 116 15 1.58e-16
c1110 101 1 1.327e-15
c1111 3 0 1.827e-15
c1112 137 136 6.36e-16
c1113 360 261 1.6e-16
c1114 1 181 4.533e-15
c1115 14 7 4.73e-16
c1116 70 417 1.58e-16
c1117 0 238 4.006e-15
c1118 159 0 3.756e-15
c1119 150 75 6.62e-16
c1120 440 4 1.58e-16
c1121 306 406 3.66e-16
c1122 184 185 2.02e-16
c1123 113 115 3.15e-16
c1124 441 1 8.3e-16
c1125 0 271 6.354e-15
c1126 1 282 3.724e-15
c1127 1 10 8.06e-16
c1128 0 511 8.06e-16
c1129 183 161 1.042e-15
c1130 51 0 8.06e-16
c1131 481 403 1.58e-16
c1132 225 247 3.15e-16
c1133 14 0 3.471e-15
c1134 498 490 3.15e-16
c1135 420 290 1.58e-16
c1136 342 397 1.58e-16
c1137 162 238 1.432e-15
c1138 357 238 1.58e-16
c1139 282 114 1.58e-16
c1140 223 15 1.275e-15
c1141 319 111 1.58e-16
c1142 0 429 3.189e-15
c1143 225 319 1.58e-16
c1144 98 182 1.58e-16
c1145 256 235 3.15e-16
c1146 493 491 1.042e-15
c1147 282 207 1.58e-16
c1148 295 167 1.58e-16
c1149 1 471 3.083e-15
c1150 98 173 4.73e-16
c1151 73 71 1.926e-15
c1152 1 263 3.083e-15
c1153 418 46 1.58e-16
c1154 0 267 3.724e-15
c1155 1 247 3.888e-15
c1156 96 83 1.58e-16
c1157 342 250 1.58e-16
c1158 1 39 1.862e-15
c1159 319 48 3.15e-16
c1160 1 395 1.862e-15
c1161 282 44 1.58e-16
c1162 342 326 1.58e-16
c1163 110 1 3.724e-15
c1164 182 180 7.96e-16
c1165 332 417 1.58e-16
c1166 510 0 5.051e-15
c1167 353 0 8.3e-16
c1168 151 139 1.58e-16
c1169 269 285 1.58e-16
c1170 0 142 3.154e-15
c1171 15 107 1.58e-16
c1172 57 0 8.3e-16
c1173 418 1 8.3e-16
c1174 381 287 6.17e-16
c1175 46 16 9.74e-16
c1176 3 48 1.275e-15
c1177 330 294 3.15e-16
c1178 245 0 8.06e-16
c1179 3 102 3.15e-16
c1180 418 144 1.9e-16
c1181 98 184 1.58e-16
c1182 269 1 8.3e-16
c1183 294 223 1.58e-16
c1184 109 133 7.5e-16
c1185 382 377 7.96e-16
c1186 1 464 6.289e-15
c1187 384 395 1.58e-16
c1188 363 380 1.58e-16
c1189 175 319 1.58e-16
c1190 290 291 8.89e-16
c1191 418 57 1.58e-16
c1192 181 182 9.74e-16
c1193 392 378 7.32e-16
c1194 0 421 8.06e-16
c1195 154 64 6.62e-16
c1196 181 173 1.58e-16
c1197 350 351 1.042e-15
c1198 367 274 1.6e-16
c1199 83 238 1.58e-16
c1200 342 311 1.58e-16
c1201 87 1 5.001e-15
c1202 90 53 9.88e-16
c1203 89 94 4.11e-16
c1204 177 0 8.06e-16
c1205 192 193 1.132e-15
c1206 413 1 1.301e-15
c1207 392 478 3.15e-16
c1208 1 16 3.724e-15
c1209 227 0 8.3e-16
c1210 285 298 3.15e-16
c1211 182 242 1.58e-16
c1212 418 19 1.58e-16
c1213 344 353 1.58e-16
c1214 424 247 2.848e-15
c1215 19 121 1.58e-16
c1216 1 379 8.06e-16
c1217 420 464 1.58e-16
c1218 432 403 1.58e-16
c1219 127 121 6.36e-16
c1220 192 367 4.8e-16
c1221 290 471 3.137e-15
c1222 1 298 9.645e-15
c1223 0 57 1.827e-15
c1224 464 384 4.48e-16
c1225 417 1 8.3e-16
c1226 96 221 1.58e-16
c1227 348 409 8.89e-16
c1228 0 145 3.756e-15
c1229 300 46 3.15e-16
c1230 124 214 1.58e-16
c1231 348 1 3.7e-15
c1232 390 1 1.327e-15
c1233 450 459 1.58e-16
c1234 59 58 3.306e-15
c1235 198 203 1.58e-16
c1236 151 299 1.58e-16
c1237 347 344 3.54e-16
c1238 81 78 1.58e-16
c1239 181 184 1.58e-16
c1240 234 263 9.54e-16
c1241 67 1 3.163e-15
c1242 92 68 9.54e-16
c1243 81 0 1.05e-15
c1244 193 197 3.15e-16
c1245 358 0 1.862e-15
c1246 158 35 3.63e-16
c1247 125 0 5.159e-15
c1248 295 0 8.3e-16
c1249 250 0 2.476e-15
c1250 305 249 1.926e-15
c1251 300 1 8.3e-16
c1252 293 297 4.6e-16
c1253 1 388 8.06e-16
c1254 1 316 3.724e-15
c1255 290 464 3.15e-16
c1256 300 144 3.15e-16
c1257 318 348 1.432e-15
c1258 324 377 1.063e-15
c1259 174 163 7.96e-16
c1260 169 0 1.444e-15
c1261 0 167 5.056e-15
c1262 269 373 5.05e-16
c1263 256 247 1.58e-16
c1264 342 0 1.327e-15
c1265 324 378 4.73e-16
c1266 0 435 3.189e-15
c1267 158 164 1.58e-16
c1268 124 1 3.289e-15
c1269 339 338 4.8e-16
c1270 206 0 8.3e-16
c1271 201 1 8.3e-16
c1272 76 77 1.6e-16
c1273 417 1 8.3e-16
c1274 217 19 3.15e-16
c1275 163 1 8.3e-16
c1276 7 106 1.263e-15
c1277 162 309 1.263e-15
c1278 443 445 9.96e-16
c1279 256 319 1.58e-16
c1280 420 316 3.15e-16
c1281 145 30 1.58e-16
c1282 282 116 1.58e-16
c1283 109 149 1.58e-16
c1284 418 167 1.58e-16
c1285 37 36 1.88e-15
c1286 342 418 1.58e-16
c1287 400 1 1.565e-15
c1288 358 0 8.3e-16
c1289 479 403 1.58e-16
c1290 1 440 3.724e-15
c1291 0 441 3.756e-15
c1292 40 39 7.32e-16
c1293 205 207 1.042e-15
c1294 1 85 7.053e-15
c1295 416 0 1.862e-15
c1296 519 510 1.132e-15
c1297 320 299 3.15e-16
c1298 144 85 1.58e-16
c1299 226 27 1.58e-16
c1300 295 0 8.3e-16
c1301 294 193 3.15e-16
c1302 96 151 1.58e-16
c1303 28 145 4.73e-16
c1304 151 226 3.15e-16
c1305 163 55 1.58e-16
c1306 57 85 1.58e-16
c1307 330 282 3.15e-16
c1308 0 37 3.756e-15
c1309 202 119 3.306e-15
c1310 290 1 1.327e-15
c1311 342 0 8.3e-16
c1312 295 113 1.58e-16
c1313 282 223 1.58e-16
c1314 7 26 1.926e-15
c1315 487 424 1.58e-16
c1316 488 486 1.58e-16
c1317 0 478 2.912e-15
c1318 169 0 1.05e-15
c1319 100 1 2.565e-15
c1320 98 97 7.96e-16
c1321 0 302 2.661e-15
c1322 158 15 1.58e-16
c1323 431 429 1.042e-15
c1324 436 435 1.042e-15
c1325 89 87 3.63e-16
c1326 125 28 8.3e-16
c1327 397 404 5.48e-16
c1328 150 0 2.893e-15
c1329 1 291 3.163e-15
c1330 0 13 8.06e-16
c1331 1 5 4.761e-15
c1332 75 85 3.15e-16
c1333 0 339 1.327e-15
c1334 256 298 2.06e-16
c1335 0 376 8.06e-16
c1336 256 390 1.58e-16
c1337 357 478 3.47e-16
c1338 275 274 1.578e-15
c1339 329 0 8.06e-16
c1340 282 107 1.58e-16
c1341 295 30 1.58e-16
c1342 304 1 1.327e-15
c1343 397 1 7.826e-15
c1344 135 226 1.88e-16
c1345 319 203 1.58e-16
c1346 300 167 1.58e-16
c1347 65 158 4.75e-16
c1348 326 404 4.6e-16
c1349 192 1 2.565e-15
c1350 96 320 1.58e-16
c1351 206 283 1.58e-16
c1352 162 307 2.5e-16
c1353 357 339 1.58e-16
c1354 64 39 1.58e-16
c1355 366 368 3.137e-15
c1356 411 347 7.32e-16
c1357 1 112 8.06e-16
c1358 295 48 1.58e-16
c1359 320 226 1.58e-16
c1360 1 237 4.616e-15
c1361 1 364 8.316e-15
c1362 96 62 3.15e-16
c1363 72 68 1.58e-16
c1364 198 195 1.96e-16
c1365 296 1 8.06e-16
c1366 285 326 1.82e-16
c1367 115 203 8.66e-16
c1368 441 283 1.58e-16
c1370 1 250 1.862e-15
c1371 193 4 1.58e-16
c1372 418 0 8.3e-16
c1373 336 417 1.063e-15
c1374 378 281 1.58e-16
c1375 219 287 3.15e-16
c1376 326 1 1.862e-15
c1377 432 387 3.15e-16
c1378 1 501 8.06e-16
c1379 1 35 5.536e-15
c1380 1 365 8.06e-16
c1381 403 394 1.58e-16
c1382 316 496 6.36e-16
c1383 0 36 3.306e-15
c1384 1 197 5.319e-15
c1385 0 119 2.6e-15
c1386 359 86 3.306e-15
c1387 7 0 4.948e-15
c1388 459 373 1.58e-16
c1389 100 358 3.15e-16
c1390 475 0 1.327e-15
c1391 492 1 3.293e-15
c1392 158 34 1.58e-16
c1393 439 417 7.96e-16
c1394 158 53 4.73e-16
c1395 175 250 1.58e-16
c1396 1 15 8.3e-16
c1397 238 320 1.58e-16
c1398 1 352 3.724e-15
c1399 89 85 1.58e-16
c1400 164 1 4.761e-15
c1401 76 1 1.327e-15
c1402 424 397 3.15e-16
c1403 283 110 1.58e-16
c1404 179 185 2.6e-16
c1406 306 238 1.58e-16
c1407 353 157 1.58e-16
c1408 311 1 8.3e-16
c1409 339 434 7.96e-16
c1410 1 371 3.548e-15
c1411 352 114 1.58e-16
c1412 24 116 6.06e-16
c1413 418 0 8.3e-16
c1414 0 113 1.444e-15
c1415 292 291 1.926e-15
c1416 449 450 2.69e-15
c1417 299 46 1.58e-16
c1418 0 121 5.051e-15
c1419 342 286 3.15e-16
c1420 1 199 1.565e-15
c1421 249 320 1.58e-16
c1422 76 55 8.3e-16
c1423 0 469 5.159e-15
c1424 120 0 8.06e-16
c1425 217 0 3.189e-15
c1426 248 229 7.96e-16
c1427 418 113 1.58e-16
c1428 270 268 1.042e-15
c1429 0 261 2.476e-15
c1430 78 87 3.15e-16
c1431 119 0 2.476e-15
c1432 113 121 4.73e-16
c1433 76 75 2.6e-16
c1434 300 0 8.3e-16
c1435 294 1 8.3e-16
c1436 1 185 3.189e-15
c1437 316 1 1.327e-15
c1438 0 337 5.076e-15
c1439 15 1 8.3e-16
c1440 129 0 3.189e-15
c1441 299 1 8.3e-16
c1442 96 143 1.58e-16
c1443 313 0 1.892e-15
c1444 171 114 4.48e-16
c1445 20 0 3.306e-15
c1446 240 242 3.15e-16
c1447 124 223 1.58e-16
c1448 322 0 8.06e-16
c1449 357 417 1.58e-16
c1450 363 366 3.15e-16
c1451 54 0 8.06e-16
c1452 299 144 3.15e-16
c1453 225 0 1.612e-15
c1454 256 397 3.15e-16
c1455 216 0 8.06e-16
c1456 405 324 9.74e-16
c1457 397 381 2.848e-15
c1458 60 46 4.6e-16
c1459 70 242 1.58e-16
c1460 169 86 8.89e-16
c1461 301 1 8.06e-16
c1462 201 1 8.3e-16
c1463 285 0 1.05e-15
c1464 313 418 1.58e-16
c1465 1 12 2.026e-15
c1466 353 58 1.58e-16
c1467 98 179 1.58e-16
c1468 318 1 3.189e-15
c1469 311 424 1.58e-16
c1470 0 470 8.06e-16
c1471 225 418 3.15e-16
c1472 403 324 9.74e-16
c1473 455 462 3.306e-15
c1474 0 262 8.06e-16
c1475 260 0 2.476e-15
c1476 395 364 1.58e-16
c1477 219 319 1.58e-16
c1478 440 1 8.3e-16
c1479 256 250 1.58e-16
c1480 319 195 3.15e-16
c1481 293 288 4.73e-16
c1482 413 414 1.58e-16
c1483 65 1 3.289e-15
c1484 173 352 3.15e-16
c1485 256 326 1.58e-16
c1486 290 330 1.58e-16
c1487 432 369 4.73e-16
c1488 209 115 7.96e-16
c1489 24 23 6.17e-16
c1490 167 170 1.58e-16
c1491 1 60 3.815e-15
c1492 124 107 8.3e-16
c1493 96 46 3.15e-16
c1494 284 282 1.926e-15
c1495 502 1 5.051e-15
c1496 48 121 1.58e-16
c1497 130 107 3.137e-15
c1498 0 313 2.6e-15
c1499 226 46 1.58e-16
c1500 294 1 8.3e-16
c1501 300 0 8.3e-16
c1502 151 140 1.58e-16
c1503 0 404 3.194e-15
c1504 1 418 4.761e-15
c1505 219 269 3.15e-16
c1506 185 1 1.862e-15
c1507 44 8 3.15e-16
c1508 418 28 4.73e-16
c1509 201 12 3.15e-16
c1510 332 389 1.132e-15
c1511 15 56 6.62e-16
c1512 225 0 3.689e-15
c1513 397 473 6.36e-16
c1514 1 493 4.591e-15
c1515 113 217 3.15e-16
c1516 330 291 3.15e-16
c1517 12 44 1.58e-16
c1518 119 48 1.58e-16
c1519 100 0 8.3e-16
c1520 98 1 8.3e-16
c1521 175 0 1.827e-15
c1522 324 274 1.58e-16
c1523 201 440 1.58e-16
c1524 151 441 1.58e-16
c1525 285 0 8.3e-16
c1526 300 113 1.58e-16
c1527 440 12 1.58e-16
c1528 0 403 1.827e-15
c1529 1 481 3.163e-15
c1530 163 78 1.58e-16
c1531 83 417 1.58e-16
c1532 96 1 1.301e-15
c1533 420 502 4.73e-16
c1534 210 19 7.32e-16
c1535 440 44 1.58e-16
c1536 506 397 6.79e-16
c1537 163 0 3.306e-15
c1538 352 184 1.58e-16
c1539 226 1 8.3e-16
c1540 96 144 1.58e-16
c1541 369 332 8.57e-16
c1542 1 173 5.151e-15
c1543 420 493 3.15e-16
c1544 78 85 2.848e-15
c1545 95 94 6.36e-16
c1546 1 315 3.163e-15
c1547 226 144 1.58e-16
c1548 34 1 7.053e-15
c1549 234 185 1.58e-16
c1550 96 57 1.58e-16
c1551 219 298 3.15e-16
c1552 0 85 1.05e-15
c1553 235 149 1.58e-16
c1554 57 226 3.34e-16
c1555 132 1 4.427e-15
c1556 292 1 8.06e-16
c1557 316 315 7.32e-16
c1558 420 481 3.15e-16
c1559 0 491 2.893e-15
c1560 469 466 3.54e-16
c1561 464 463 7.96e-16
c1562 96 55 3.15e-16
c1563 306 309 1.58e-16
c1564 300 30 1.58e-16
c1565 295 203 1.58e-16
c1566 255 179 6.62e-16
c1567 299 167 1.58e-16
c1568 450 447 2.848e-15
c1569 109 157 1.58e-16
c1570 271 268 6.36e-16
c1571 96 75 1.58e-16
c1572 181 1 8.3e-16
c1573 98 1 2.565e-15
c1574 100 0 8.3e-16
c1575 260 261 3.54e-16
c1576 363 441 1.58e-16
c1577 300 48 1.58e-16
c1578 255 257 1.042e-15
c1579 86 0 2.6e-15
c1580 393 378 1.926e-15
c1581 282 1 8.3e-16
c1582 1 242 5.854e-15
c1583 24 118 7.96e-16
c1584 363 377 9.74e-16
c1585 366 267 1.58e-16
c1586 0 507 8.06e-16
c1587 424 0 1.327e-15
c1588 369 275 1.58e-16
c1589 1 70 4.109e-15
c1590 470 466 4.8e-16
c1591 243 1 8.06e-16
c1592 139 0 2.144e-15
c1593 132 1 1.862e-15
c1594 441 104 1.58e-16
c1595 100 261 1.58e-16
c1596 256 0 8.3e-16
c1597 1 406 5.854e-15
c1598 162 237 7.32e-16
c1599 432 1 8.3e-16
c1600 458 0 1.327e-15
c1601 293 287 3.15e-16
c1602 109 319 1.58e-16
c1603 341 344 6.62e-16
c1604 0 373 1.892e-15
c1605 1 260 3.289e-15
c1606 440 364 1.204e-15
c1607 446 445 7.96e-16
c1608 448 395 6.36e-16
c1609 64 164 1.82e-16
c1610 86 87 1.03e-16
c1611 420 70 3.15e-16
c1612 173 182 1.58e-16
c1613 256 418 1.58e-16
c1614 0 444 8.06e-16
c1615 181 1 2.565e-15
c1616 62 39 1.58e-16
c1617 57 249 3.15e-16
c1618 116 114 3.15e-16
c1619 411 344 4.73e-16
c1620 96 167 4.73e-16
c1621 282 1 8.3e-16
c1622 157 149 1.58e-16
c1623 330 1 2.565e-15
c1624 96 342 1.58e-16
c1625 226 167 1.58e-16
c1626 175 163 9.74e-16
c1627 227 145 1.58e-16
c1628 111 5 1.58e-16
c1629 1 223 1.862e-15
c1630 306 307 8.89e-16
c1631 432 384 3.15e-16
c1632 429 427 2.848e-15
c1633 170 78 3.15e-16
c1634 1 332 2.514e-15
c1635 397 414 3.15e-16
c1636 256 0 8.3e-16
c1637 100 1 8.3e-16
c1638 170 0 3.154e-15
c1639 488 487 1.58e-16
c1640 1 477 1.565e-15
c1641 381 0 5.056e-15
c1642 139 0 1.05e-15
c1643 222 1 8.06e-16
c1644 250 251 1.6e-16
c1645 82 71 7.96e-16
c1646 184 182 1.58e-16
c1647 234 181 1.58e-16
c1648 498 397 3.15e-16
c1649 166 1 4.616e-15
c1650 76 78 5.11e-16
c1651 173 184 3.15e-16
c1652 0 455 4.492e-15
c1653 154 75 1.042e-15
c1654 299 0 8.3e-16
c1655 83 164 3.15e-16
c1656 72 53 3.15e-16
c1657 417 27 1.58e-16
c1658 76 0 2.6e-15
c1659 308 1 8.06e-16
c1660 420 332 3.98e-16
c1661 151 417 1.58e-16
c1662 304 407 3.15e-16
c1663 432 290 1.58e-16
c1664 490 500 1.58e-16
c1665 1 479 3.163e-15
c1666 342 238 1.58e-16
c1667 151 362 1.58e-16
c1668 269 372 3.15e-16
c1669 287 288 1.658e-15
c1670 311 494 3.306e-15
c1671 460 386 3.306e-15
c1672 418 25 1.58e-16
c1673 1 190 8.06e-16
c1674 350 352 6.36e-16
c1675 256 300 1.58e-16
c1676 219 295 1.58e-16
c1677 441 267 1.58e-16
c1678 269 265 3.15e-16
c1679 1 380 3.815e-15
c1680 437 411 3.6e-16
c1681 392 369 7.09e-16
c1682 210 0 3.719e-15
c1683 109 142 1.58e-16
c1684 1 275 3.293e-15
c1685 86 85 1.96e-16
c1686 219 326 1.58e-16
c1687 420 479 3.15e-16
c1688 283 15 1.58e-16
c1689 268 167 6.62e-16
c1690 334 231 7.96e-16
c1691 299 0 8.3e-16
c1692 319 0 8.3e-16
c1693 218 217 1.042e-15
c1694 244 169 1.926e-15
c1695 0 147 8.06e-16
c1696 432 304 3.15e-16
c1697 133 145 3.15e-16
c1698 0 58 6.319e-15
c1699 96 0 8.3e-16
c1700 432 395 3.15e-16
c1701 299 113 1.58e-16
c1702 124 1 8.3e-16
c1703 100 86 2.6e-16
c1704 0 200 2.893e-15
c1705 226 0 3.306e-15
c1706 417 320 3.15e-16
c1707 363 362 7.32e-16
c1708 447 373 3.15e-16
c1709 98 0 1.862e-15
c1710 3 0 1.892e-15
c1711 159 0 8.3e-16
c1712 1 462 1.565e-15
c1713 247 303 1.58e-16
c1714 306 417 1.58e-16
c1715 352 240 1.58e-16
c1716 83 65 1.58e-16
c1717 441 1 8.3e-16
c1718 385 0 2.912e-15
c1719 64 53 1.58e-16
c1720 141 1 8.06e-16
c1721 109 145 6.3e-16
c1722 39 46 1.58e-16
c1723 283 294 1.58e-16
c1724 70 352 1.58e-16
c1725 192 368 6.36e-16
c1726 249 302 1.275e-15
c1727 299 30 1.58e-16
c1728 293 298 1.58e-16
c1729 155 226 3.15e-16
c1730 300 203 1.58e-16
c1731 39 61 1.58e-16
c1732 96 78 3.15e-16
c1733 0 105 2.144e-15
c1734 238 0 3.756e-15
c1735 352 158 1.58e-16
c1736 24 1 1.862e-15
c1737 96 0 8.3e-16
c1738 201 193 1.58e-16
c1739 299 48 1.58e-16
c1740 12 193 3.15e-16
c1741 39 1 7.684e-15
c1742 124 1 1.327e-15
c1743 0 186 1.05e-15
c1744 226 0 8.3e-16
c1745 130 1 3.083e-15
c1746 193 44 1.58e-16
c1747 14 119 6.73e-16
c1748 144 39 1.58e-16
c1749 110 1 8.3e-16
c1750 415 1 1.301e-15
c1751 440 193 3.15e-16
c1752 0 353 4.006e-15
c1753 151 274 3.15e-16
c1754 464 332 1.58e-16
c1755 70 1 2.247e-15
c1756 418 414 3.15e-16
c1757 1 505 5.854e-15
c1758 502 513 6.36e-16
c1759 1 187 1.565e-15
c1760 57 39 5.74e-16
c1761 164 27 1.58e-16
c1762 113 226 1.58e-16
c1763 316 70 1.58e-16
c1764 1 392 3.724e-15
c1765 0 369 5.617e-15
c1766 249 0 1.327e-15
c1767 86 170 1.58e-16
c1768 151 192 1.58e-16
c1769 39 55 4.73e-16
c1770 219 0 8.3e-16
c1771 70 114 1.58e-16
c1772 347 0 2.6e-15
c1773 311 488 1.58e-16
c1774 0 414 3.719e-15
c1775 395 275 1.58e-16
c1776 109 295 1.58e-16
c1777 432 316 1.58e-16
c1778 420 505 3.15e-16
c1779 1 277 4.59e-15
c1780 75 39 1.74e-16
c1781 162 242 1.58e-16
c1782 284 1 8.06e-16
c1783 105 0 1.05e-15
c1784 352 179 3.15e-16
c1785 7 145 1.58e-16
c1786 347 418 1.58e-16
c1787 420 392 3.15e-16
c1788 357 369 3.15e-16
c1789 208 115 3.306e-15
c1790 140 167 3.15e-16
c1791 158 114 3.39e-16
c1792 283 4 1.58e-16
c1793 225 226 7.32e-16
c1794 312 309 1.926e-15
c1795 288 379 1.926e-15
c1796 0 428 2.893e-15
c1797 226 30 1.58e-16
c1798 109 169 1.275e-15
c1799 418 227 1.9e-16
c1800 298 288 6.3e-16
c1801 227 121 1.58e-16
c1802 332 1 2.565e-15
c1803 62 35 1.58e-16
c1804 145 0 8.3e-16
c1805 231 1 3.724e-15
c1806 386 387 8.89e-16
c1807 119 195 1.03e-16
c1808 219 0 8.3e-16
c1809 96 1 8.3e-16
c1810 487 486 2.848e-15
c1811 347 0 1.892e-15
c1812 155 154 6.36e-16
c1813 214 1 5.854e-15
c1814 345 1 1.565e-15
c1815 339 435 9.74e-16
c1816 437 413 3.15e-16
c1817 363 192 3.15e-16
c1818 226 28 1.58e-16
c1819 490 397 2.78e-16
c1820 159 161 1.58e-16
c1821 81 0 1.862e-15
c1822 352 1 8.3e-16
c1823 399 386 6.36e-16
c1825 320 164 1.58e-16
c1826 1 239 8.06e-16
c1827 240 182 9.74e-16
c1828 86 84 6.36e-16
c1829 281 282 8.89e-16
c1830 492 493 2.69e-15
c1831 68 1 5.051e-15
c1832 154 0 2.893e-15
c1833 227 129 1.58e-16
c1834 417 46 1.58e-16
c1835 0 297 2.912e-15
c1836 164 62 1.58e-16
c1837 136 0 2.893e-15
c1838 319 235 3.15e-16
c1839 342 378 1.58e-16
c1840 70 182 1.58e-16
c1841 225 238 3.15e-16
c1842 70 173 1.58e-16
c1843 282 283 1.88e-15
c1844 437 390 3.66e-16
c1845 70 315 1.421e-15
c1846 397 468 6.69e-16
c1847 250 149 6.73e-16
c1848 219 217 2.69e-15
c1849 48 105 1.58e-16
c1850 376 377 7.96e-16
c1851 417 1 8.3e-16
c1852 124 126 1.6e-16
c1853 7 295 1.58e-16
c1854 219 300 1.58e-16
c1855 151 294 1.58e-16
c1856 256 299 1.58e-16
c1857 1 238 1.301e-15
c1858 342 339 1.58e-16
c1859 417 144 1.58e-16
c1860 173 158 9.74e-16
c1861 275 1 4.109e-15
c1862 217 227 3.15e-16
c1863 259 182 7.96e-16
c1864 225 249 1.58e-16
c1865 437 487 3.15e-16
c1866 57 417 1.58e-16
c1867 352 1 8.3e-16
c1868 320 15 1.58e-16
c1869 70 184 1.58e-16
c1870 441 188 1.58e-16
c1871 353 85 1.58e-16
c1872 295 0 8.3e-16
c1873 293 295 3.15e-16
c1874 413 411 8.3e-16
c1875 418 133 1.58e-16
c1876 357 348 1.58e-16
c1877 1 207 4.591e-15
c1878 417 19 1.9e-16
c1879 175 238 6.17e-16
c1880 293 326 1.58e-16
c1881 50 15 1.58e-16
c1882 140 0 1.862e-15
c1883 201 1 3.293e-15
c1884 206 0 1.327e-15
c1885 501 70 1.926e-15
c1886 101 0 1.827e-15
c1887 12 1 1.862e-15
c1888 109 0 1.612e-15
c1889 96 86 1.58e-16
c1890 420 0 8.3e-16
c1891 357 1 8.3e-16
c1892 290 324 1.58e-16
c1893 455 363 8.89e-16
c1894 440 1 8.3e-16
c1895 441 0 8.3e-16
c1896 0 384 4.006e-15
c1897 179 182 7.75e-16
c1898 234 352 1.58e-16
c1899 171 1 3.163e-15
c1900 173 179 1.289e-15
c1901 418 109 1.58e-16
c1902 392 464 1.58e-16
c1903 486 397 3.15e-16
c1904 109 121 1.58e-16
c1905 278 113 1.926e-15
c1906 0 94 3.189e-15
c1907 189 193 4.6e-16
c1908 182 257 1.132e-15
c1909 287 298 1.58e-16
c1910 424 238 1.58e-16
c1911 275 323 7.96e-16
c1912 369 386 1.58e-16
c1913 267 274 6.73e-16
c1914 1 366 3.163e-15
c1915 256 96 6.62e-16
c1916 357 420 1.58e-16
c1917 1 398 3.083e-15
c1918 96 381 3.15e-16
c1919 225 423 6.62e-16
c1920 1 114 1.023e-14
c1921 41 40 1.88e-15
c1922 397 288 1.58e-16
c1923 299 203 1.58e-16
c1924 50 294 1.58e-16
c1925 274 271 1.58e-16
c1926 495 311 7.96e-16
c1927 35 46 3.15e-16
c1928 294 104 1.58e-16
c1929 192 267 9.32e-16
c1930 0 290 4.545e-15
c1931 140 0 3.754e-15
c1932 184 179 1.58e-16
c1933 1 182 4.427e-15
c1934 101 0 1.892e-15
c1935 12 1 8.3e-16
c1936 1 234 1.862e-15
c1937 81 161 1.58e-16
c1938 68 89 8.3e-16
c1939 173 1 2.691e-15
c1940 1 44 1.862e-15
c1941 247 319 2.38e-16
c1942 288 295 1.58e-16
c1943 151 132 3.15e-16
c1944 440 1 8.3e-16
c1945 441 0 8.3e-16
c1946 0 265 3.154e-15
c1947 140 113 4.6e-16
c1948 206 113 3.15e-16
c1949 417 167 1.58e-16
c1950 1 83 4.376e-15
c1951 49 0 8.06e-16
c1952 342 417 1.58e-16
c1953 164 46 1.58e-16
c1954 326 288 4.73e-16
c1955 62 53 1.58e-16
c1956 35 1 1.327e-15
c1957 437 397 1.58e-16
c1958 490 503 3.15e-16
c1959 144 35 3.47e-16
c1960 256 238 1.58e-16
c1961 313 408 1.03e-16
c1962 225 309 1.58e-16
c1963 311 486 3.15e-16
c1964 137 214 3.15e-16
c1965 319 115 1.58e-16
c1966 222 221 1.926e-15
c1967 455 454 1.03e-16
c1968 1 466 7.098e-15
c1969 39 78 3.15e-16
c1970 1 184 9.066e-15
c1971 0 372 3.154e-15
c1972 1 427 8.29e-15
c1973 109 300 1.58e-16
c1974 420 83 3.15e-16
c1975 319 3 3.15e-16
c1976 0 39 1.444e-15
c1977 164 1 8.3e-16
c1978 0 395 2.6e-15
c1979 293 0 5.298e-15
c1980 437 326 1.58e-16
c1981 110 0 3.306e-15
c1982 182 1 1.862e-15
c1983 286 297 1.58e-16
c1984 519 1 4.591e-15
c1985 173 1 4.427e-15
c1986 226 25 1.58e-16
c1987 132 135 6.06e-16
c1988 256 249 1.58e-16
c1989 206 285 1.58e-16
c1990 1 408 5.001e-15
c1991 74 46 7.96e-16
c1992 441 111 1.58e-16
c1993 57 164 1.58e-16
c1994 20 49 7.96e-16
c1995 357 304 1.58e-16
c1996 0 496 2.893e-15
c1997 122 1 3.083e-15
c1998 7 119 3.54e-16
c1999 418 0 8.3e-16
c2000 15 46 4.03e-16
c2001 132 320 1.58e-16
c2002 204 48 1.926e-15
c2003 310 0 3.194e-15
c2004 336 1 4.427e-15
c2005 285 441 1.58e-16
c2006 206 1 8.3e-16
c2007 139 227 1.58e-16
c2008 164 55 3.15e-16
c2009 0 464 5.051e-15
c2010 412 1 8.06e-16
c2011 441 48 1.58e-16
c2012 447 445 1.289e-15
c2013 420 519 3.15e-16
c2014 411 397 3.15e-16
c2015 153 76 3.306e-15
c2016 234 182 1.58e-16
c2017 1 386 1.862e-15
c2018 441 1 8.3e-16
c2019 75 164 1.58e-16
c2020 234 173 3.15e-16
c2021 0 344 5.051e-15
c2022 415 414 1.58e-16
c2023 437 311 1.58e-16
c2024 87 0 2.912e-15
c2025 184 1 3.293e-15
c2026 0 303 3.154e-15
c2027 324 1 2.565e-15
c2028 293 0 1.862e-15
c2029 416 1 5.854e-15
c2030 0 16 3.306e-15
c2031 15 1 8.316e-15
c2032 285 378 3.15e-16
c2033 15 144 1.58e-16
c2034 339 337 3.54e-16
c2035 275 330 3.15e-16
c2036 1 377 5.051e-15
c2037 357 464 1.58e-16
c2038 369 363 1.59e-15
c2039 110 111 2.038e-15
c2040 313 307 7.32e-16
c2041 336 318 1.58e-16
c2042 418 344 4.73e-16
c2043 397 287 1.58e-16
c2044 223 1 4.427e-15
c2045 1 378 5.677e-15
c2046 417 0 8.3e-16
c2047 225 307 1.263e-15
c2048 162 352 3.15e-16
c2049 386 384 4.18e-16
c2050 0 194 8.06e-16
c2051 7 300 1.58e-16
c2052 162 239 1.926e-15
c2053 219 299 1.58e-16
c2054 282 104 3.15e-16
c2055 516 397 5.05e-16
c2056 234 184 1.9e-16
c2057 261 263 3.137e-15
c2058 15 55 3.15e-16
c2059 288 0 5.116e-15
c2060 348 343 1.58e-16
c2061 67 0 2.493e-15
c2062 116 1 5.677e-15
c2063 1 189 3.841e-15
c2064 19 15 1.58e-16
c2065 92 90 3.137e-15
c2066 78 68 1.58e-16
c2067 65 1 1.327e-15
c2068 128 0 8.06e-16
c2069 274 167 3.15e-16
c2070 326 287 1.58e-16
c2071 339 1 1.862e-15
c2072 1 229 3.163e-15
c2073 390 298 7.32e-16
c2074 300 0 8.3e-16
c2075 294 1 8.3e-16
c2076 0 316 4.462e-15
c2077 510 506 9.74e-16
c2078 31 32 2.038e-15
c2079 70 240 1.125e-15
c2080 432 407 3.15e-16
c2081 223 224 1.926e-15
c2082 466 471 6.36e-16
c2083 1 211 8.06e-16
c2084 34 46 1.58e-16
c2085 53 46 1.58e-16
c2086 246 0 8.06e-16
c2087 290 386 1.58e-16
c2088 252 184 6.36e-16
c2089 162 1 5.536e-15
c2090 357 1 3.293e-15
c2091 40 42 1.926e-15
c2092 65 55 1.58e-16
c2093 201 0 8.3e-16
c2094 151 1 8.3e-16
c2095 417 0 8.3e-16
c2096 163 0 8.3e-16
c2097 357 316 1.58e-16
c2098 0 288 4.127e-15
c2099 96 353 1.58e-16
c2100 82 0 8.06e-16
c2101 61 53 1.58e-16
c2102 432 70 1.58e-16
c2103 294 19 1.58e-16
c2104 401 0 8.06e-16
c2105 479 481 3.15e-16
c2106 0 440 3.306e-15
c2107 34 1 1.301e-15
c2108 0 85 6.15e-15
c2109 1 53 1.1439e-14
c2110 417 113 1.58e-16
c2111 83 352 1.58e-16
c2112 34 144 1.58e-16
c2113 144 53 3.15e-16
c2114 109 139 1.58e-16
c2115 464 466 9.74e-16
c2116 357 318 3.15e-16
c2117 64 114 1.58e-16
c2118 1 107 5.051e-15
c2119 57 53 1.9e-16
c2120 397 247 3.15e-16
c2121 200 195 6.62e-16
c2122 167 15 1.58e-16
c2123 437 0 1.327e-15
c2124 96 227 3.15e-16
c2125 281 1 1.327e-15
c2126 341 0 2.893e-15
c2127 100 0 1.327e-15
c2128 98 1 1.862e-15
c2129 386 395 3.15e-16
c2130 226 227 2.038e-15
c2131 55 53 4.73e-16
c2132 313 417 1.58e-16
c2133 500 397 3.15e-16
c2134 1 363 1.862e-15
c2135 225 417 1.58e-16
c2136 1 193 5.151e-15
c2137 417 30 1.58e-16
c2138 192 188 1.58e-16
c2139 1 283 4.761e-15
c2140 83 1 3.289e-15
c2141 293 286 1.58e-16
c2142 0 5 3.756e-15
c2143 1 4 3.724e-15
c2144 75 53 3.15e-16
c2145 0 513 2.893e-15
c2146 256 378 1.58e-16
c2147 432 332 2.46e-16
c2148 319 295 4.73e-16
c2149 151 290 1.58e-16
c2150 316 83 1.58e-16
c2151 256 478 3.15e-16
c2152 250 319 1.58e-16
c2153 1 306 3.289e-15
c2154 411 418 3.15e-16
c2155 0 47 8.06e-16
c2156 83 114 1.9e-16
c2157 305 1 8.06e-16
c2158 1 417 3.724e-15
c2159 287 0 2.771e-15
c2160 417 28 1.58e-16
c2161 142 145 3.15e-16
c2162 295 115 1.58e-16
c2163 221 214 1.58e-16
c2164 294 167 1.58e-16
c2165 162 173 1.58e-16
c2166 363 384 1.58e-16
c2167 109 299 1.58e-16
c2168 192 0 1.327e-15
c2169 201 283 1.58e-16
c2170 151 291 1.58e-16
c2171 1 362 4.616e-15
c2172 413 397 6.3e-16
c2173 283 12 1.58e-16
c2174 0 237 3.719e-15
c2175 1 240 3.163e-15
c2176 0 364 5.581e-15
c2177 71 68 1.58e-16
c2178 283 44 1.58e-16
c2179 420 306 1.58e-16
c2180 440 283 1.58e-16
c2181 411 0 4.043e-15
c2183 70 1 8.3e-16
c2184 50 24 1.58e-16
c2185 311 247 1.58e-16
c2186 282 1 8.3e-16
c2187 24 104 1.132e-15
c2188 132 19 1.58e-16
c2189 124 50 1.58e-16
c2190 502 505 3.15e-16
c2191 193 1 8.3e-16
c2192 342 387 1.58e-16
c2193 397 390 3.15e-16
c2194 0 35 3.439e-15
c2195 324 330 1.58e-16
c2196 162 184 1.58e-16
c2197 287 0 3.689e-15
c2198 0 197 3.189e-15
c2199 355 0 8.06e-16
c2200 492 0 1.327e-15
c2201 497 1 3.293e-15
c2202 98 358 1.132e-15
c2203 163 161 3.15e-16
c2204 173 178 7.96e-16
c2205 288 286 1.58e-16
c2206 1 454 5.001e-15
c2207 0 463 8.06e-16
c2208 326 298 6.3e-16
c2209 0 15 8.3e-16
c2210 193 191 7.96e-16
c2211 89 53 3.15e-16
c2212 164 0 3.756e-15
c2213 76 0 2.476e-15
c2214 213 50 7.96e-16
c2215 269 371 1.46e-16
c2216 487 397 3.15e-16
c2217 179 257 1.58e-16
c2219 83 173 1.58e-16
c2220 488 238 1.58e-16
c2221 517 502 6.36e-16
c2222 405 1 5.854e-15
c2223 125 145 3.15e-16
c2224 411 436 6.36e-16
c2225 96 109 1.58e-16
c2226 70 1 8.3e-16
c2227 151 214 1.58e-16
c2228 231 1 1.327e-15
c2229 109 226 1.58e-16
c2230 403 1 2.565e-15
c2231 151 352 1.58e-16
c2232 7 299 2.14e-16
c2233 288 380 1.58e-16
c2234 326 487 3.15e-16
c2235 220 1 1.565e-15
c2236 247 0 8.3e-16
c2237 100 161 1.58e-16
c2238 363 395 1.66e-16
c2239 1 179 6.214e-15
c2240 0 360 8.06e-16
c2241 68 95 3.137e-15
c2242 158 1 3.724e-15
c2243 294 0 8.3e-16
c2244 83 184 1.58e-16
c2245 306 304 1.58e-16
c2246 84 0 2.893e-15
c2247 0 185 4.492e-15
c2248 1 257 4.591e-15
c2249 0 319 3.306e-15
c2250 1 343 5.319e-15
c2251 285 274 1.58e-16
c2252 428 427 1.042e-15
c2253 15 0 8.3e-16
c2254 299 0 8.3e-16
c2255 70 234 1.58e-16
c2256 418 247 1.58e-16
c2257 132 131 7.96e-16
c2258 256 417 2.06e-16
c2259 474 476 1.042e-15
c2260 478 482 7.96e-16
c2261 164 30 1.58e-16
c2262 1 274 1.327e-15
c2263 469 381 3.15e-16
c2264 1 480 5.854e-15
c2265 418 319 1.58e-16
c2266 503 500 3.47e-16
c2267 285 192 1.58e-16
c2268 113 15 1.58e-16
c2269 269 0 1.327e-15
c2270 151 1 8.3e-16
c2271 428 408 6.62e-16
c2272 0 3 1.862e-15
c2273 339 340 6.36e-16
c2274 311 487 2.06e-16
c2275 135 214 3.15e-16
c2276 282 167 1.58e-16
c2277 455 450 2.02e-16
c2278 1 192 7.047e-15
c2279 0 247 3.724e-15
c2280 432 505 3.15e-16
c2281 164 28 1.58e-16
c2282 65 78 1.58e-16
c2283 136 133 6.62e-16
c2284 115 121 1.58e-16
c2285 320 214 1.58e-16
c2286 319 119 1.58e-16
c2287 0 448 2.893e-15
c2288 416 414 3.15e-16
c2289 65 0 1.827e-15
c2290 420 480 3.15e-16
c2291 432 392 1.58e-16
c2292 342 369 1.58e-16
c2293 0 60 3.194e-15
c2294 179 1 2.565e-15
c2295 24 46 3.15e-16
c2296 502 0 7.092e-15
c2297 281 330 1.58e-16
c2298 14 110 3.15e-16
c2299 294 0 8.3e-16
c2300 352 62 1.58e-16
c2301 185 0 2.6e-15
c2302 50 214 1.132e-15
c2303 469 473 3.137e-15
c2304 0 493 3.189e-15
c2305 1 146 8.06e-16
c2306 266 101 3.306e-15
c2307 298 0 1.892e-15
c2308 15 30 2.22e-16
c2309 330 283 3.15e-16
c2310 197 48 3.15e-16
c2311 98 0 8.3e-16
c2312 151 440 1.58e-16
c2313 219 441 1.58e-16
c2314 269 0 8.3e-16
c2315 170 161 3.15e-16
c2316 294 113 1.58e-16
c2317 140 227 3.15e-16
c2318 283 223 1.58e-16
c2319 287 286 7.32e-16
c2320 0 481 2.912e-15
c2321 224 1 8.06e-16
c2322 24 1 3.189e-15
c2323 335 319 7.96e-16
c2324 96 0 1.05e-15
c2325 48 15 3.15e-16
c2326 418 298 3.15e-16
c2327 43 30 7.96e-16
c2328 234 179 1.58e-16
c2329 226 0 8.3e-16
c2330 24 144 3.15e-16
c2331 392 332 1.58e-16
c2332 353 39 1.58e-16
c2333 417 25 1.58e-16
c2334 78 53 4.73e-16
c2335 1 320 4.761e-15
c2336 15 28 3.79e-16
c2337 413 0 1.05e-15
c2338 326 397 3.15e-16
c2339 392 477 3.306e-15
c2340 34 0 6.15e-15
c2341 270 1 4.591e-15
c2342 132 0 3.189e-15
c2343 319 300 4.73e-16
c2344 173 230 7.32e-16
c2345 306 1 1.327e-15
c2346 348 435 1.58e-16
c2347 402 324 7.96e-16
c2348 0 298 6.494e-15
c2349 294 111 1.58e-16
c2350 320 114 1.58e-16
c2351 24 19 3.15e-16
c2352 347 346 6.36e-16
c2353 124 19 7.82e-16
c2354 390 0 1.892e-15
c2355 62 114 1.58e-16
c2356 300 115 1.58e-16
c2357 457 384 6.62e-16
c2358 461 447 1.042e-15
c2359 151 173 3.15e-16
c2360 181 0 8.3e-16
c2361 234 1 3.189e-15
c2362 98 0 1.327e-15
c2363 363 440 1.58e-16
c2364 294 48 3.15e-16
c2365 50 114 1.58e-16
c2366 311 397 4.73e-16
c2367 282 0 8.3e-16
c2368 1 358 2.565e-15
c2369 0 242 3.154e-15
c2370 397 396 4.8e-16
c2371 370 267 9.74e-16
c2372 502 83 1.58e-16
c2373 0 180 8.06e-16
c2374 104 12 1.74e-16
c2375 342 348 3.15e-16
c2376 0 70 3.055e-15
c2377 41 1 4.761e-15
c2378 132 0 1.862e-15
c2379 440 104 1.58e-16
c2380 151 364 1.58e-16
c2381 252 1 3.083e-15
c2382 255 0 2.893e-15
c2383 298 300 1.58e-16
c2384 324 332 3.15e-16
c2385 1 387 3.163e-15
c2386 420 358 1.58e-16
c2387 432 0 8.3e-16
c2388 342 1 8.3e-16
c2389 418 145 1.58e-16
c2390 220 137 3.306e-15
c2391 159 85 3.31e-16
c2392 132 113 1.58e-16
c2393 70 162 4.73e-16
c2394 357 70 1.58e-16
c2395 28 34 7.63e-16
c2396 392 483 7.96e-16
c2397 181 0 1.327e-15
c2398 0 99 8.06e-16
c2399 486 238 3.15e-16
c2400 319 5 1.58e-16
c2401 411 415 5.11e-16
c2402 282 0 8.3e-16
c2403 283 193 4.11e-16
c2404 109 140 1.58e-16
c2405 124 167 1.58e-16
c2406 206 109 1.58e-16
c2407 96 437 1.58e-16
c2408 357 432 1.58e-16
c2409 352 46 1.58e-16
c2410 111 4 1.58e-16
c2411 417 414 1.047e-15
c2412 129 145 3.15e-16
c2413 269 447 4.73e-16
c2414 342 384 3.15e-16
c2415 293 398 9.54e-16
c2416 410 1 8.06e-16
c2417 0 332 2.144e-15
c2418 98 1 8.3e-16
c2419 282 113 1.58e-16
c2420 137 1 3.189e-15
c2421 267 1 1.301e-15
c2422 363 364 1.263e-15
c2423 419 1 8.06e-16
c2424 316 429 1.58e-16
c2425 64 158 1.58e-16
c2426 261 181 5.11e-16
c2427 125 129 5.11e-16
c2428 166 0 3.719e-15
c2429 503 397 3.47e-16
c2430 275 324 9.74e-16
c2431 151 330 3.15e-16
c2432 397 418 3.15e-16
c2433 487 406 3.15e-16
c2434 71 53 3.15e-16
c2435 352 1 8.3e-16
c2436 1 271 5.051e-15
c2437 0 295 3.756e-15
c2438 0 11 8.06e-16
c2439 86 185 1.58e-16
c2440 151 223 1.58e-16
c2441 250 0 8.3e-16
c2442 357 332 1.58e-16
c2443 219 417 1.58e-16
c2444 390 476 1.58e-16
c2445 164 25 1.58e-16
c2446 326 0 1.327e-15
c2447 347 417 1.58e-16
c2448 0 375 8.06e-16
c2449 342 290 1.58e-16
c2450 83 70 3.15e-16
c2451 0 479 3.649e-15
c2452 248 0 8.06e-16
c2453 230 229 1.58e-16
c2454 298 286 4.73e-16
c2455 219 362 1.58e-16
c2456 437 238 1.58e-16
c2457 295 121 1.58e-16
c2458 282 111 3.15e-16
c2459 250 418 1.58e-16
c2460 417 227 3.47e-16
c2461 109 110 8.89e-16
c2462 397 0 3.189e-15
c2463 19 214 4.03e-16
c2464 0 472 8.06e-16
c2465 326 418 3.15e-16
c2466 352 55 1.58e-16
c2467 453 373 3.306e-15
c2468 440 267 1.58e-16
c2469 206 265 1.58e-16
c2470 1 389 5.854e-15
c2471 1 108 8.06e-16
c2472 282 48 1.58e-16
c2473 83 158 1.58e-16
c2474 0 275 1.327e-15
c2475 137 1 1.862e-15
c2476 235 236 1.926e-15
c2478 372 377 1.132e-15
c2479 0 250 2.6e-15
c2480 152 1 5.319e-15
c2481 50 116 1.58e-16
c2482 311 0 1.892e-15
c2483 185 183 6.36e-16
c2484 104 116 1.58e-16
c2485 398 288 3.137e-15
c2486 342 304 1.58e-16
c2487 369 1 6.062e-15
c2488 326 0 1.862e-15
c2489 256 387 3.15e-16
c2490 76 58 4.73e-16
c2491 57 1 8.3e-16
c2492 145 85 1.58e-16
c2493 0 205 2.893e-15
c2494 1 8 3.724e-15
c2495 158 172 7.96e-16
c2496 203 15 1.58e-16
c2497 81 163 3.15e-16
c2498 173 143 1.275e-15
c2499 162 1 4.109e-15
c2500 342 395 3.15e-16
c2501 320 223 3.15e-16
c2502 144 114 1.58e-16
c2503 124 0 8.3e-16
c2504 311 418 1.58e-16
c2505 0 483 8.06e-16
c2506 228 1 8.06e-16
c2507 12 1 2.565e-15
c2508 238 235 3.15e-16
c2509 399 381 1.042e-15
c2510 57 114 1.9e-16
c2511 81 85 1.58e-16
c2512 175 242 1.132e-15
c2513 1 450 5.319e-15
c2514 44 1 2.565e-15
c2515 324 394 8.97e-16
c2516 95 53 9.54e-16
c2517 87 94 3.15e-16
c2518 441 0 8.3e-16
c2519 440 1 8.3e-16
c2521 319 299 4.73e-16
c2522 295 300 4.73e-16
c2523 309 303 1.58e-16
c2524 19 114 1.58e-16
c2525 311 0 8.3e-16
c2526 511 411 1.6e-16
c2527 0 371 2.661e-15
c2528 397 406 3.47e-16
c2529 143 184 1.58e-16
c2530 213 0 8.06e-16
c2531 0 396 8.06e-16
c2532 1 42 8.06e-16
c2533 75 114 3.15e-16
c2534 435 409 1.58e-16
c2535 432 386 4.73e-16
c2536 352 167 1.58e-16
c2537 7 110 3.15e-16
c2538 293 378 1.82e-16
c2539 294 203 6.3e-16
c2540 299 115 1.58e-16
c2541 447 459 1.58e-16
c2542 450 384 1.58e-16
c2543 485 479 6.36e-16
c2544 24 0 1.862e-15
c2545 162 1 1.327e-15
c2546 50 107 1.58e-16
c2547 39 0 7.799e-15
c2548 124 0 2.476e-15
c2549 93 90 1.6e-16
c2550 91 89 1.6e-16
c2551 31 1 3.724e-15
c2552 358 1 2.026e-15
c2553 283 1 8.3e-16
c2554 83 1 8.3e-16
c2555 353 164 1.58e-16
c2556 110 0 8.3e-16
c2557 326 406 9.74e-16
c2558 219 274 1.58e-16
c2559 64 1 3.7e-15
c2560 413 415 3.15e-16
c2561 0 505 3.154e-15
c2562 510 411 5.11e-16
c2563 417 109 1.58e-16
c2564 124 113 1.58e-16
c2565 418 0 8.3e-16
c2566 369 373 1.58e-16
c2567 397 476 3.79e-16
c2568 351 353 1.58e-16
c2569 100 397 3.15e-16
c2570 0 392 4.462e-15
c2571 1 167 7.515e-15
c2572 219 192 1.58e-16
c2573 298 299 8.89e-16
c2574 162 234 1.58e-16
c2575 342 1 3.293e-15
c2576 1 348 3.163e-15
c2577 48 190 1.926e-15
c2578 247 226 9.74e-16
c2579 289 1 8.06e-16
c2580 493 306 1.58e-16
c2581 285 1 8.3e-16
c2582 418 121 1.74e-16
c2583 86 166 1.58e-16
c2584 346 344 1.042e-15
c2585 96 319 1.58e-16
c2586 342 316 1.58e-16
c2587 227 164 1.58e-16
c2588 167 114 6.17e-16
c2589 312 1 8.06e-16
c2590 120 121 4.8e-16
c2591 24 111 1.58e-16
c2592 357 392 1.58e-16
c2593 256 369 6.17e-16
c2594 94 85 1.58e-16
c2595 24 30 3.15e-16
c2596 96 58 4.73e-16
c2597 385 399 6.62e-16
c2598 517 0 2.893e-15
c2599 510 516 9.21e-16
c2600 369 381 3.15e-16
c2601 119 121 5.11e-16
c2602 288 377 7.32e-16
c2603 283 1 8.3e-16
c2604 83 1 8.3e-16
c2605 327 0 8.06e-16
c2606 0 418 3.756e-15
c2607 342 318 3.15e-16
c2608 326 286 3.15e-16
c2609 378 288 1.58e-16
c2610 120 119 1.6e-16
c2611 24 48 1.132e-15
c2612 96 159 1.58e-16
c2613 335 0 8.06e-16
c2614 330 271 3.15e-16
c2615 197 195 2.848e-15
c2616 420 1 1.301e-15
c2617 247 238 1.58e-16
c2618 221 1 3.163e-15
c2619 214 0 3.154e-15
c2620 104 193 1.58e-16
c2621 384 1 2.565e-15
c2622 231 230 3.15e-16
c2623 1 302 3.548e-15
c2624 130 28 9.54e-16
c2625 352 0 8.3e-16
c2626 319 105 1.58e-16
c2627 238 319 1.58e-16
c2628 90 1 3.189e-15
c2629 68 0 6.437e-15
c2630 227 15 1.58e-16
c2631 83 234 1.58e-16
c2632 0 300 3.756e-15
c2633 358 173 3.15e-16
c2634 186 185 2.6e-16
c2635 96 298 3.15e-16
c2636 217 121 3.15e-16
c2637 357 336 1.58e-16
c2638 437 478 3.15e-16
c2639 505 83 1.289e-15
c2640 70 320 1.58e-16
c2641 469 468 3.54e-16
c2642 1 424 3.289e-15
c2643 418 300 1.58e-16
c2644 247 249 1.58e-16
c2645 431 250 6.36e-16
c2646 300 121 1.58e-16
c2647 1 272 1.565e-15
c2648 116 19 1.432e-15
c2649 173 167 1.58e-16
c2650 290 1 8.3e-16
c2651 282 203 1.58e-16
c2652 39 79 3.137e-15
c2653 417 0 8.3e-16
c2654 293 417 1.58e-16
c2655 249 319 1.58e-16
c2656 219 294 1.58e-16
c2657 437 339 1.58e-16
c2658 357 324 1.58e-16
c2659 352 155 1.58e-16
c2660 260 0 8.3e-16
c2661 411 412 1.926e-15
c2662 294 195 3.15e-16
c2663 12 188 1.58e-16
c2664 1 373 5.151e-15
c2665 91 78 4.8e-16
c2666 432 306 1.74e-16
c2667 420 424 1.58e-16
c2668 158 62 1.58e-16
c2670 225 304 4.18e-16
c2671 352 0 8.3e-16
c2672 1 230 4.616e-15
c2673 152 64 1.58e-16
c2674 440 188 1.58e-16
c2675 0 436 2.893e-15
c2676 353 53 1.58e-16
c2678 0 207 3.189e-15
c2679 1 23 3.815e-15
c2680 201 0 1.327e-15
c2681 151 1 8.3e-16
c2682 151 275 3.15e-16
c2683 12 0 1.862e-15
c2684 417 344 4.73e-16
c2685 98 186 3.15e-16
c2686 100 0 1.862e-15
c2687 0 406 3.154e-15
c2688 1 304 5.151e-15
c2689 231 320 1.58e-16
c2690 384 373 3.15e-16
c2691 357 0 8.3e-16
c2692 256 1 8.3e-16
c2693 358 356 1.042e-15
c2694 415 397 4.73e-16
c2695 1 381 2.514e-15
c2696 76 150 6.36e-16
c2697 440 0 8.3e-16
c2698 1 395 1.327e-15
c2699 0 260 1.827e-15
c2700 0 286 3.719e-15
c2701 324 281 1.58e-16
c2702 423 247 1.042e-15
c2703 87 85 3.15e-16
c2704 171 0 2.912e-15
c2705 100 418 3.15e-16
c2706 269 366 3.15e-16
c2707 480 481 1.132e-15
c2708 96 145 1.58e-16
c2709 287 378 1.58e-16
c2710 487 238 3.15e-16
c2711 413 510 4.73e-16
c2712 416 516 9.74e-16
c2713 517 519 1.042e-15
c2714 19 107 1.58e-16
c2715 295 299 1.58e-16
c2716 226 145 1.58e-16
c2717 411 339 1.58e-16
c2718 19 23 1.58e-16
c2719 127 107 9.54e-16
c2720 1 370 5.854e-15
c2721 19 211 1.926e-15
c2722 256 420 1.58e-16
c2723 14 282 3.15e-16
c2724 1 113 1.862e-15
c2725 96 81 1.58e-16
c2726 326 422 7.96e-16
c2727 0 114 7.16e-15
c2728 381 384 1.58e-16
c2729 100 0 8.3e-16
c2730 35 36 7.32e-16
c2731 168 1 8.06e-16
c2732 427 247 9.74e-16
c2733 1 473 3.083e-15
c2734 109 15 1.58e-16
c2735 135 1 6.214e-15
c2736 151 1 3.293e-15
c2737 363 275 7.82e-16
c2738 12 0 8.3e-16
c2739 0 182 3.189e-15
c2740 1 261 1.327e-15
c2741 70 429 1.58e-16
c2742 90 89 5.11e-16
c2743 173 0 2.273e-15
c2744 0 44 1.444e-15
c2745 320 1 8.3e-16
c2746 192 265 1.58e-16
c2747 424 304 2.02e-16
c2748 113 207 1.58e-16
c2749 223 167 1.578e-15
c2750 440 0 8.3e-16
c2751 0 279 6.18e-15
c2752 1 337 3.189e-15
c2753 313 1 1.327e-15
c2754 1 506 3.163e-15
c2755 0 83 4.006e-15
c2756 193 1 8.3e-16
c2757 432 429 3.005e-15
c2758 35 0 1.892e-15
c2759 225 1 2.247e-15
c2760 437 469 1.58e-16
c2761 96 397 1.58e-16
c2762 132 227 1.58e-16
c2763 50 1 4.376e-15
c2764 353 242 1.58e-16
c2765 290 381 3.15e-16
c2766 0 485 2.893e-15
c2767 430 313 3.306e-15
c2768 285 1 1.301e-15
c2769 175 352 1.58e-16
c2770 137 221 8.89e-16
c2771 0 466 3.189e-15
c2772 0 184 3.724e-15
c2773 163 85 3.15e-16
c2774 260 262 1.6e-16
c2775 109 294 1.58e-16
c2776 83 162 1.58e-16
c2777 0 380 3.194e-15
c2778 1 409 7.541e-15
c2779 395 373 1.58e-16
c2780 452 364 6.62e-16
c2781 357 83 1.58e-16
c2782 420 506 3.15e-16
c2783 111 8 3.15e-16
c2784 173 155 3.63e-16
c2785 318 337 3.54e-16
c2786 17 46 1.58e-16
c2787 34 133 3.15e-16
c2788 164 0 8.3e-16
c2789 135 1 2.565e-15
c2790 96 326 1.58e-16
c2791 182 0 1.862e-15
c2792 205 203 6.62e-16
c2793 231 143 7.32e-16
c2794 24 25 1.58e-16
c2795 12 111 1.58e-16
c2796 441 319 1.58e-16
c2797 519 0 3.189e-15
c2798 316 1 8.3e-16
c2799 48 114 1.58e-16
c2800 173 0 3.189e-15
c2801 333 231 7.96e-16
c2802 1 430 1.565e-15
c2803 0 431 2.893e-15
c2804 320 1 8.3e-16
c2805 158 46 1.58e-16
c2806 111 44 1.58e-16
c2807 124 203 1.58e-16
c2808 325 0 8.06e-16
c2809 201 285 1.58e-16
c2810 206 269 4.73e-16
c2811 44 30 1.132e-15
c2812 440 111 1.58e-16
c2813 70 1 1.327e-15
c2814 473 290 9.54e-16
c2815 1 62 1.301e-15
c2816 101 3 2.6e-16
c2817 28 114 4.73e-16
c2818 12 48 1.58e-16
c2819 397 238 4.73e-16
c2820 53 37 1.58e-16
c2821 1 17 4.761e-15
c2822 100 260 1.58e-16
c2823 175 1 3.289e-15
c2824 285 440 1.58e-16
c2825 201 1 8.3e-16
c2826 269 441 6.3e-16
c2827 50 1 3.289e-15
c2828 109 34 1.58e-16
c2829 7 15 1.58e-16
c2830 441 3 3.15e-16
c2831 318 1 4.495e-15
c2832 381 395 3.18e-16
c2833 109 53 3.15e-16
c2834 44 102 1.432e-15
c2835 104 1 5.854e-15
c2836 440 48 2.38e-16
c2837 349 1 1.565e-15
c2838 450 364 1.58e-16
c2839 158 1 8.3e-16
c2840 440 1 8.3e-16
c2841 0 386 2.6e-15
c2842 66 53 1.926e-15
c2843 74 0 8.06e-16
c2844 86 352 3.15e-16
c2845 261 173 6.73e-16
c2846 281 283 1.58e-16
c2847 184 0 1.327e-15
c2848 0 299 3.306e-15
c2849 250 238 1.58e-16
c2850 1 18 8.06e-16
c2851 15 0 5.581e-15
c2852 344 351 2.848e-15
c2853 416 413 7.63e-16
c2854 57 158 1.58e-16
c2855 256 464 1.58e-16
c2856 437 403 1.58e-16
c2857 464 381 6.06e-16
c2858 469 287 6.73e-16
c2859 1 494 1.565e-15
c2860 223 0 2.771e-15
c2861 143 1 8.218e-15
c2862 418 299 3.66e-16
c2863 0 43 8.06e-16
c2864 299 121 1.58e-16
c2865 151 137 3.15e-16
c2866 158 55 4.73e-16
c2867 159 39 1.58e-16
c2868 256 352 1.58e-16
c2869 151 152 2.69e-15
c2870 151 324 1.58e-16
c2871 480 479 1.58e-16
c2872 140 142 9.74e-16
c2873 0 189 4.036e-15
c2874 28 31 9.74e-16
c2875 75 158 1.58e-16
c2876 116 0 4.637e-15
c2877 86 1 1.862e-15
c2878 14 24 4.73e-16
c2879 84 87 6.62e-16
c2880 65 0 1.892e-15
c2881 287 383 7.96e-16
c2882 378 298 1.905e-15
c2883 275 271 1.58e-16
c2884 415 0 1.05e-15
c2885 0 422 8.06e-16
c2886 0 229 2.912e-15
c2887 397 398 6.36e-16
c2888 311 238 8.66e-16
c2889 294 0 8.3e-16
c2890 293 294 1.289e-15
c2891 1 498 4.591e-15
c2892 413 339 3.005e-15
c2893 176 114 7.96e-16
c2894 478 390 1.58e-16
c2895 86 114 1.58e-16
c2896 223 155 7.32e-16
c2897 347 348 1.03e-16
c2898 53 36 1.132e-15
c2899 144 146 1.926e-15
c2900 504 503 1.926e-15
c2901 170 85 3.15e-16
c2902 256 1 8.3e-16
c2903 96 0 8.3e-16
c2904 143 1 1.327e-15
c2905 175 173 1.58e-16
c2906 151 0 8.3e-16
c2907 219 1 8.3e-16
c2908 135 137 1.03e-16
c2909 336 320 1.58e-16
c2910 70 167 1.58e-16
c2911 1 364 2.247e-15
c2912 109 282 1.58e-16
c2913 420 498 3.15e-16
c2914 342 70 1.58e-16
c2915 76 85 1.58e-16
c2916 164 161 3.15e-16
c2917 96 418 1.58e-16
c2918 142 39 1.58e-16
c2919 34 0 1.05e-15
c2920 0 53 8.322e-15
c2921 418 226 1.74e-16
c2922 116 111 1.58e-16
c2923 521 510 7.96e-16
c2924 226 121 1.58e-16
c2925 300 299 2.207e-15
c2926 245 140 7.96e-16
c2927 342 432 1.58e-16
c2928 214 203 1.58e-16
c2929 57 1 8.3e-16
c2930 188 193 1.58e-16
c2931 219 124 1.58e-16
c2932 234 143 1.58e-16
c2933 109 166 7.32e-16
c2934 417 247 1.58e-16
c2935 8 9 1.892e-15
c2936 0 107 6.437e-15
c2937 116 48 1.58e-16
c2938 175 184 1.58e-16
c2939 397 427 4.73e-16
c2940 200 119 6.36e-16
c2941 96 0 8.3e-16
c2942 19 1 4.109e-15
c2943 417 319 1.58e-16
c2944 238 0 1.612e-15
c2945 98 0 1.862e-15
c2946 505 429 3.15e-16
c2947 450 448 1.042e-15
c2948 226 129 1.58e-16
c2949 113 107 1.58e-16
c2950 86 182 1.58e-16
c2951 0 363 1.444e-15
c2953 86 173 1.58e-16
c2954 288 294 8.89e-16
c2955 285 330 3.15e-16
c2956 397 408 4.39e-16
c2957 0 193 3.689e-15
c2958 92 1 3.083e-15
c2959 84 85 1.042e-15
c2960 250 427 1.03e-16
c2961 0 4 3.306e-15
c2962 342 332 3.15e-16
c2963 418 238 1.58e-16
c2964 241 185 7.32e-16
c2965 143 252 3.137e-15
c2966 145 39 1.58e-16
c2967 1 330 1.862e-15
c2968 1 144 3.724e-15
c2969 1 488 5.001e-15
c2970 0 306 1.827e-15
c2971 151 281 1.58e-16
c2972 269 362 3.15e-16
c2973 1 391 8.06e-16
c2974 0 268 2.893e-15
c2975 249 0 1.444e-15
c2976 57 1 8.3e-16
c2977 256 182 1.58e-16
c2978 217 226 3.15e-16
c2979 111 107 3.15e-16
c2980 56 46 1.042e-15
c2981 189 48 7.32e-16
c2982 162 320 1.58e-16
c2983 96 300 1.58e-16
c2984 151 283 3.15e-16
c2985 364 373 1.03e-16
c2986 7 282 3.15e-16
c2987 0 238 1.05e-15
c2988 416 397 4.73e-16
c2989 86 184 1.58e-16
c2990 0 240 2.912e-15
c2991 1 445 6.452e-15
c2992 19 1 2.247e-15
c2993 65 161 1.58e-16
c2994 357 306 1.58e-16
c2995 420 488 3.15e-16
c2996 127 1 3.083e-15
c2997 207 203 1.58e-16
c2998 298 417 1.58e-16
c2999 48 107 1.58e-16
c3000 70 0 8.3e-16
c3001 48 23 1.58e-16
c3002 75 1 5.726e-15
c3003 282 0 8.3e-16
c3004 193 0 8.3e-16
c3005 397 478 3.47e-16
c3006 437 387 3.15e-16
c3007 96 163 1.58e-16
c3008 1 167 2.247e-15
c3009 340 1 3.083e-15
c3010 275 167 1.58e-16
c3011 311 309 7.32e-16
c3012 498 496 1.042e-15
c3013 118 0 8.06e-16
c3014 1 202 1.565e-15
c3015 356 86 6.36e-16
c3016 96 85 3.15e-16
c3017 497 0 1.327e-15
c3018 518 1 3.293e-15
c3019 339 397 3.15e-16
c3020 259 0 8.06e-16
c3021 0 454 2.912e-15
c3022 198 199 3.306e-15
c3023 352 353 1.193e-15
c3024 83 320 1.58e-16
c3025 318 340 3.137e-15
c3026 373 330 7.32e-16
c3027 70 78 1.58e-16
c3028 31 25 7.32e-16
c3029 212 294 1.58e-16
c3030 0 366 3.733e-15
c3031 109 24 4.73e-16
c3032 70 0 8.3e-16
c3033 321 319 1.926e-15
c3034 1 32 4.761e-15
c3035 151 221 3.15e-16
c3036 231 0 1.892e-15
c3037 193 111 1.58e-16
c3038 96 286 3.15e-16
c3039 167 1 4.761e-15
c3040 14 8 9.74e-16
c3041 283 104 1.58e-16
c3042 128 125 1.6e-16
c3043 98 161 1.58e-16
c3044 0 179 4.006e-15
c3045 186 1 1.301e-15
c3046 158 0 3.306e-15
c3047 193 48 3.15e-16
c3048 417 145 1.58e-16
c3049 123 0 8.06e-16
c3050 421 324 7.96e-16
c3051 0 423 2.893e-15
c3052 14 44 3.15e-16
c3053 1 188 5.001e-15
c3054 0 257 3.189e-15
c3055 72 1 4.761e-15
c3056 0 309 4.637e-15
c3057 1 353 6.214e-15
c3058 256 223 4.73e-16
c3059 1 490 1.2276e-14
c3060 0 509 8.06e-16
c3061 40 1 3.724e-15
c3062 498 316 1.171e-15
c3063 311 307 1.58e-16
c3064 0 480 3.154e-15
c3065 269 192 4.73e-16
c3066 353 114 1.58e-16
c3067 206 0 8.3e-16
c3068 219 1 8.3e-16
c3069 324 57 1.58e-16
c3070 1 407 3.815e-15
c3071 159 164 1.58e-16
c3072 243 241 1.926e-15
c3073 1 266 1.565e-15
c3074 0 101 2.6e-15
c3075 347 1 1.862e-15
c3076 493 424 1.58e-16
c3077 137 19 1.58e-16
c3078 363 386 1.58e-16
c3079 455 461 6.36e-16
c3080 1 468 4.616e-15
c3081 395 445 1.58e-16
c3082 111 17 3.15e-16
c3083 0 427 5.051e-15
c3084 420 490 7.88e-16
c3085 17 30 3.15e-16
c3086 441 0 8.3e-16
c3087 319 197 3.15e-16
c3088 1 443 3.815e-15
c3089 40 55 9.74e-16
c3090 51 31 7.96e-16
c3091 29 1 8.06e-16
c3092 437 369 5.21e-16
c3093 179 0 1.327e-15
c3094 152 75 2.848e-15
c3095 319 15 1.58e-16
c3096 70 1 8.3e-16
c3097 24 7 1.362e-15
c3098 96 139 1.58e-16
c3099 0 408 2.912e-15
c3100 397 417 3.15e-16
c3101 420 468 3.15e-16
c3102 469 397 1.58e-16
c3103 227 114 1.58e-16
c3104 139 226 1.58e-16
c3105 264 3 6.62e-16
c3106 347 318 3.15e-16
c3107 416 418 1.58e-16
c3108 142 35 1.58e-16
c3109 15 58 1.03e-16
c3110 122 14 9.54e-16
c3111 12 195 9.74e-16
c3112 165 163 1.926e-15
c3113 115 15 1.58e-16
c3114 212 132 9.74e-16
c3115 96 76 1.58e-16
c3116 219 440 1.58e-16
c3117 206 0 8.3e-16
c3118 432 1 3.293e-15
c3119 175 240 6.17e-16
c3120 348 344 1.58e-16
c3121 103 44 1.926e-15
c3122 155 1 1.327e-15
c3123 346 0 2.893e-15
c3124 24 0 3.754e-15
c3125 425 304 3.306e-15
c3126 450 275 1.58e-16
c3127 69 1 8.06e-16
c3128 158 28 1.58e-16
c3129 250 417 1.58e-16
c3130 418 378 4.73e-16
c3131 166 161 3.15e-16
c3132 0 441 8.3e-16
c3133 0 457 2.893e-15
c3134 345 337 3.306e-15
c3135 225 231 1.58e-16
c3136 68 94 1.58e-16
c3137 1 297 3.163e-15
c3138 0 307 4.215e-15
c3139 339 0 1.862e-15
c3140 416 0 3.154e-15
c3141 369 474 6.62e-16
c3142 138 1 1.565e-15
c3143 353 182 1.58e-16
c3144 64 1 1.301e-15
c3145 357 57 1.58e-16
c3146 173 353 1.58e-16
c3147 515 416 7.96e-16
c3148 319 294 4.73e-16
c3149 70 71 7.32e-16
c3150 342 336 1.58e-16
c3151 0 377 5.616e-15
c3152 320 230 3.15e-16
c3153 464 465 7.96e-16
c3154 290 468 6.73e-16
c3155 1 486 6.582e-15
c3156 113 1 8.3e-16
c3157 251 184 4.8e-16
c3158 339 418 1.58e-16
c3159 0 378 4.637e-15
c3160 1 332 5.151e-15
c3161 117 116 1.926e-15
c3162 151 135 3.15e-16
c3163 151 363 1.58e-16
c3164 320 27 1.58e-16
c3165 35 145 3.15e-16
c3166 294 115 3.15e-16
c3167 65 159 3.15e-16
c3168 109 352 1.58e-16
c3169 0 191 8.06e-16
c3170 151 320 1.58e-16
c3171 96 299 1.58e-16
c3172 342 324 1.58e-16
c3173 293 290 1.58e-16
c3174 294 3 3.15e-16
c3175 186 184 1.58e-16
c3176 261 1 1.862e-15
c3177 234 0 3.754e-15
c3178 287 282 9.74e-16
c3179 311 417 4.7e-16
c3180 78 92 6.36e-16
c3181 155 1 1.862e-15
c3182 14 116 3.15e-16
c3183 420 486 3.15e-16
c3184 432 424 1.58e-16
c3185 353 184 1.58e-16
c3186 339 0 1.862e-15
c3187 369 287 4.19e-16
c3188 0 358 1.327e-15
c3189 75 64 1.58e-16
c3190 151 50 1.58e-16
c3191 283 1 8.3e-16
c3192 293 291 3.15e-16
c3193 83 1 2.565e-15
c3194 413 512 9.54e-16
c3195 225 1 1.327e-15
c3196 397 403 7.05e-16
c3197 133 114 3.15e-16
c3198 41 0 3.756e-15
c3199 490 496 6.62e-16
c3200 285 275 3.15e-16
c3201 219 364 1.58e-16
c3202 67 39 1.432e-15
c3203 109 1 2.247e-15
c3204 113 1 3.815e-15
c3205 1 48 3.724e-15
c3206 81 164 1.58e-16
c3207 96 60 5.48e-16
c3208 256 240 3.15e-16
c3209 357 358 2.848e-15
c3210 384 288 1.58e-16
c3211 342 0 8.3e-16
c3212 437 1 8.3e-16
c3213 33 31 1.926e-15
c3214 254 240 7.96e-16
c3215 159 53 4.73e-16
c3216 1 275 8.3e-16
c3217 440 445 9.74e-16
c3218 256 70 1.58e-16
c3219 293 395 6.73e-16
c3220 326 403 1.58e-16
c3221 109 114 3.15e-16
c3222 298 387 1.263e-15
c3223 319 4 1.58e-16
c3224 162 167 1.58e-16
c3225 267 368 9.54e-16
c3226 464 468 3.15e-16
c3227 256 432 1.58e-16
c3228 432 381 3.15e-16
c3229 1 38 8.06e-16
c3230 15 145 1.58e-16
c3231 96 226 3.15e-16
c3232 1 280 8.06e-16
c3233 458 459 2.69e-15
c3234 1 111 4.761e-15
c3235 8 13 7.96e-16
c3236 163 39 1.58e-16
c3237 175 1 4.376e-15
c3238 417 0 8.3e-16
c3239 290 288 1.58e-16
c3240 193 203 1.58e-16
c3241 3 4 7.32e-16
c3242 137 0 4.492e-15
c3243 143 230 1.58e-16
c3244 304 303 1.58e-16
c3245 137 138 3.306e-15
c3246 326 274 9.74e-16
c3247 360 181 4.8e-16
c3248 261 234 3.54e-16
c3249 68 87 3.15e-16
c3250 48 1 8.3e-16
c3251 128 129 4.8e-16
c3252 387 388 1.926e-15
c3253 418 417 2.049e-15
c3254 1 102 3.548e-15
c3255 417 121 1.58e-16
c3256 288 291 1.263e-15
c3257 441 5 1.58e-16
c3258 219 330 3.15e-16
c3259 91 0 8.06e-16
c3260 1 265 6.582e-15
c3261 352 0 8.3e-16
c3262 431 427 6.62e-16
c3263 28 1 7.013e-15
c3264 151 143 3.15e-16
c3265 219 223 1.58e-16
c3266 510 415 3.15e-16
c3267 1 411 1.327e-15
c3268 256 332 3.15e-16
c3269 256 231 1.58e-16
c3270 478 476 3.47e-16
c3271 142 53 3.15e-16
c3272 319 282 4.73e-16
c3273 437 290 3.15e-16
c3274 316 490 8.66e-16
c3275 378 286 3.15e-16
c3276 151 267 1.58e-16
c3277 0 417 3.306e-15
c3278 417 129 1.58e-16
c3279 256 179 1.58e-16
c3280 311 491 6.36e-16
c3281 282 115 1.58e-16
c3282 19 221 1.275e-15
c3283 283 167 1.58e-16
c3284 83 167 1.58e-16
c3285 109 173 3.15e-16
c3286 1 287 1.862e-15
c3287 455 459 3.15e-16
c3288 457 386 6.36e-16
c3289 67 68 7.32e-16
c3290 175 1 2.565e-15
c3291 445 364 3.15e-16
c3292 275 373 2.02e-16
c3293 201 265 1.58e-16
c3294 342 83 1.58e-16
c3295 0 362 3.719e-15
c3296 1 394 6.329e-15
c3297 420 411 1.58e-16
c3298 395 288 6.69e-16
c3299 86 1 1.327e-15
c3300 265 12 2.69e-15
c3301 256 257 2.848e-15
c3302 27 46 3.31e-16
c3303 0 452 2.893e-15
c3304 137 0 2.6e-15
c3305 110 5 1.58e-16
c3306 344 352 2.02e-16
c3307 293 1 8.368e-15
c3308 269 369 3.15e-16
c3309 126 0 8.06e-16
c3310 7 8 8.89e-16
c3311 516 1 8.778e-15
c3313 380 377 6.17e-16
c3314 295 15 1.58e-16
c3315 158 25 1.58e-16
c3316 152 0 3.189e-15
c3317 140 139 6.06e-16
c3318 0 383 8.06e-16
c3319 392 1 1.327e-15
c3320 1 499 1.565e-15
c3321 34 145 4.73e-16
c3322 113 137 1.58e-16
c3323 330 297 1.132e-15
c3324 7 44 1.58e-16
c3325 287 384 1.244e-15
c3326 1 27 4.616e-15
c3327 0 8 3.306e-15
c3328 175 234 1.58e-16
c3329 109 184 1.58e-16
c3330 162 0 3.055e-15
c3331 256 1 3.293e-15
c3332 310 1 3.815e-15
c3333 405 418 4.39e-16
c3334 417 300 1.58e-16
c3335 338 337 1.6e-16
c3336 420 516 4.73e-16
c3337 12 0 1.327e-15
c3338 336 337 6.73e-16
c3339 369 298 1.275e-15
c3340 0 450 3.189e-15
c3341 44 0 1.327e-15
c3342 350 353 6.62e-16
c3343 1 344 9.019e-15
c3344 68 85 3.15e-16
c3345 1 303 5.854e-15
c3346 440 0 8.3e-16
c3347 369 390 1.58e-16
c3348 86 1 8.3e-16
c3349 151 57 1.58e-16
c3351 173 149 2.06e-16
c3352 295 294 2.364e-15
c3353 437 464 1.58e-16
c3354 475 476 2.69e-15
c3355 405 0 3.154e-15
c3356 283 188 1.58e-16
c3357 397 387 3.15e-16
c3358 270 271 1.013e-15
c3359 274 0 3.306e-15
c3360 109 116 1.58e-16
c3361 151 19 1.58e-16
c3362 342 386 4.73e-16
c3363 320 46 1.9e-16
c3364 403 0 1.327e-15
c3365 336 1 3.289e-15
c3366 76 39 6.69e-16
c3367 318 344 6.3e-16
c3368 285 324 1.58e-16
c3369 162 0 1.892e-15
c3370 192 0 8.3e-16
c3371 288 1 5.822e-15
c3372 140 147 7.96e-16
c3373 155 64 1.03e-16
c3374 160 158 1.926e-15
c3375 258 185 3.306e-15
c3376 122 7 3.137e-15
c3377 86 234 1.58e-16
c3378 31 0 3.306e-15
c3379 50 46 1.58e-16
c3380 193 195 3.15e-16
c3381 283 0 8.3e-16
c3382 83 0 8.3e-16
c3383 1 324 3.724e-15
c3384 62 61 1.275e-15
c3385 0 351 3.189e-15
c3386 64 0 1.862e-15
c3387 320 1 8.3e-16
c3388 418 164 1.58e-16
c3389 416 415 3.15e-16
c3390 510 511 4.8e-16
c3391 100 417 3.15e-16
c3392 1 500 4.616e-15
c3393 62 1 2.247e-15
c3394 320 144 1.58e-16
c3395 471 287 9.54e-16
c3396 98 397 3.15e-16
c3397 1 203 1.4523e-14
c3398 70 353 1.58e-16
c3399 0 274 2.476e-15
c3400 144 62 1.58e-16
c3401 106 107 7.32e-16
c3402 57 320 1.58e-16
c3403 417 286 1.58e-16
c3404 50 1 2.565e-15
c3405 287 395 1.58e-16
c3406 0 264 2.893e-15
c3407 285 0 8.3e-16
c3408 269 1 8.3e-16
c3409 493 488 1.58e-16
c3410 57 62 1.58e-16
c3411 135 19 1.88e-16
c3412 374 330 1.926e-15
c3413 50 144 1.58e-16
c3414 22 1 8.06e-16
c3415 342 343 2.848e-15
c3416 0 192 4.006e-15
c3417 437 316 7.16e-16
c3418 0 273 3.719e-15
c3419 124 319 1.58e-16
c3420 420 500 3.15e-16
c3421 357 313 1.58e-16
c3422 171 161 6.47e-16
c3423 178 0 8.06e-16
c3424 320 19 1.58e-16
c3425 28 29 1.926e-15
c3426 0 15 1.612e-15
c3427 353 158 1.58e-16
c3428 109 107 2.62e-16
c3429 280 223 1.926e-15
c3430 71 72 2.038e-15
c3431 212 214 1.741e-15
c3432 205 115 6.36e-16
c3433 357 225 3.15e-16
c3434 94 53 3.15e-16
c3435 83 78 1.58e-16
c3436 413 1 6.401e-15
c3437 151 167 9.45e-16
c3438 339 415 3.15e-16
c3439 369 459 1.58e-16
c3440 283 0 8.3e-16
c3441 83 0 8.3e-16
c3442 464 287 1.58e-16
c3443 96 140 3.15e-16
c3444 75 62 1.58e-16
c3445 50 19 3.15e-16
c3446 418 15 1.9e-16
c3447 7 116 3.15e-16
c3448 15 121 1.58e-16
c3449 140 226 3.15e-16
c3450 269 384 3.15e-16
c3451 161 114 1.58e-16
c3452 397 389 3.15e-16
c3453 197 119 1.96e-16
c3454 357 1 8.3e-16
c3455 283 113 1.58e-16
c3456 1 390 3.289e-15
c3457 221 0 2.493e-15
c3458 98 94 9.74e-16
c3459 420 413 4.73e-16
c3460 172 0 8.06e-16
c3461 411 409 1.03e-16
c3462 90 0 5.159e-15
c3463 15 16 7.32e-16
c3464 0 294 3.306e-15
c3465 369 397 6.3e-16
c3466 96 378 1.58e-16
c3467 1 514 1.565e-15
c3468 4 6 1.926e-15
c3469 21 1 4.761e-15
c3470 317 1 8.06e-16
c3471 282 295 3.15e-16
c3472 175 162 3.15e-16
c3473 420 390 1.58e-16
c3474 1 487 3.327e-15
c3475 0 424 1.827e-15
c3476 83 313 3.15e-16
c3477 149 229 4.6e-16
c3478 328 0 8.06e-16
c3479 96 39 4.73e-16
c3480 285 281 1.58e-16
c3481 293 330 4.73e-16
c3482 283 111 1.58e-16
c3483 163 164 1.88e-15
c3484 287 1 4.427e-15
c3485 320 167 1.58e-16
c3486 386 450 1.58e-16
c3487 143 144 8.89e-16
c3488 355 352 7.96e-16
c3489 1 281 5.536e-15
c3490 256 324 1.58e-16
c3491 186 1 8.3e-16
c3492 201 198 1.58e-16
c3493 411 318 1.432e-15
c3494 117 1 8.06e-16
c3495 294 119 1.58e-16
c3496 283 48 1.58e-16
c3497 164 85 3.15e-16
c3498 0 373 4.427e-15
c3499 342 306 3.66e-16
c3500 420 487 3.15e-16
c3501 182 161 4.6e-16
c3502 352 157 1.58e-16
c3503 353 1 8.3e-16
c3504 83 1 8.3e-16
c3506 173 161 4.6e-16
c3507 0 230 3.719e-15
c3508 300 15 3.15e-16
c3509 290 298 4.7e-16
c3510 160 1 8.06e-16
c3511 218 137 6.36e-16
c3512 502 490 1.58e-16
c3514 418 34 1.58e-16
c3515 34 121 2.69e-15
c3516 14 1 5.151e-15
c3517 316 499 3.306e-15
c3518 1 46 6.452e-15
c3519 0 23 3.194e-15
c3520 151 0 8.3e-16
c3521 219 1 3.293e-15
c3522 244 1 8.06e-16
c3523 219 275 3.15e-16
c3524 269 395 3.15e-16
c3525 98 0 8.3e-16
c3526 0 387 2.493e-15
c3527 144 46 1.58e-16
c3528 1 195 8.29e-15
c3529 417 299 5.74e-16
c3530 256 0 8.3e-16
c3531 467 1 1.301e-15
c3532 83 175 1.58e-16
c3533 0 381 2.144e-15
c3534 1 459 4.591e-15
c3535 1 227 4.761e-15
c3536 57 46 2.848e-15
c3537 61 1 4.427e-15
c3538 238 307 1.421e-15
c3539 70 109 4.7e-16
c3540 426 247 7.96e-16
c3541 87 53 3.15e-16
c3542 184 161 2.69e-15
c3543 129 34 1.58e-16
c3544 399 0 2.893e-15
c3545 269 370 1.46e-16
c3546 186 1 3.7e-15
c3547 24 145 1.58e-16
c3548 0 97 8.06e-16
c3549 83 71 9.74e-16
c3550 416 510 1.58e-16
c3551 294 300 3.15e-16
c3552 288 330 4.73e-16
c3553 19 46 3.15e-16
c3554 144 1 8.3e-16
c3555 353 1 8.3e-16
c3556 256 162 1.58e-16
c3557 397 348 3.15e-16
c3558 256 357 1.58e-16
c3559 317 315 1.926e-15
c3560 331 0 8.06e-16
c3561 352 58 1.58e-16
c3562 151 155 3.15e-16
c3563 75 46 9.74e-16
c3564 57 1 3.293e-15
c3565 55 61 3.15e-16
c3566 124 125 3.54e-16
c3567 274 279 4.6e-16
c3568 459 384 1.58e-16
c3569 98 0 8.3e-16
c3570 57 144 1.58e-16
c3571 1 397 4.533e-15
c3572 479 488 2.6e-16
c3573 132 121 1.58e-16
c3574 135 0 4.006e-15
c3575 151 0 1.327e-15
c3576 247 1 8.3e-16
c3577 386 1 3.189e-15
c3578 55 1 1.023e-14
c3579 67 53 3.15e-16
c3580 0 181 1.862e-15
c3581 65 85 1.58e-16
c3582 19 1 4.616e-15
c3583 1 103 8.06e-16
c3584 320 0 8.3e-16
c3585 19 144 1.58e-16
c3586 153 1 1.565e-15
c3587 143 167 1.58e-16
c3588 88 1 1.565e-15
c3589 234 353 1.58e-16
c3590 0 282 3.306e-15
c3591 1 319 3.724e-15
c3592 227 1 8.3e-16
c3593 75 1 2.565e-15
c3594 336 340 9.54e-16
c3595 385 324 4.39e-16
c3596 510 339 1.58e-16
c3597 0 506 2.912e-15
c3598 193 0 8.3e-16
c3599 96 417 1.58e-16
c3600 96 469 1.58e-16
c3601 420 397 1.58e-16
c3602 417 226 3.15e-16
c3603 132 129 9.74e-16
c3604 50 0 4.006e-15
c3605 267 167 3.15e-16
c3606 1 368 3.083e-15
c3607 1 326 2.514e-15
c3608 490 70 1.59e-15
c3609 282 121 1.58e-16
c3610 269 1 3.293e-15
c3611 1 3 3.7e-15
c3612 493 486 3.15e-16
c3613 319 207 1.58e-16
c3614 271 167 8.78e-16
c3615 455 447 1.96e-16
c3616 163 53 1.58e-16
c3617 325 274 7.96e-16
c3618 24 295 1.58e-16
c3619 76 164 1.58e-16
c3620 0 389 3.154e-15
c3621 275 445 2.69e-15
c3622 256 83 1.58e-16
c3623 319 12 1.58e-16
c3624 100 185 4.7e-16
c3625 124 295 1.58e-16
c3626 318 319 7.32e-16
c3627 27 30 3.15e-16
c3628 1 451 1.565e-15
c3629 135 0 1.327e-15
c3630 319 44 1.58e-16
c3631 7 17 3.15e-16
c3632 207 115 1.171e-15
c3633 420 326 1.58e-16
c3634 53 85 1.236e-15
c3635 173 157 3.15e-16
c3636 440 319 1.58e-16
c3637 159 114 3.15e-16
c3638 294 5 1.58e-16
c3639 320 0 8.3e-16
c3640 132 217 9.74e-16
c3641 151 285 3.15e-16
c3642 201 269 4.73e-16
c3643 70 0 1.892e-15
c3644 1 311 3.724e-15
c3645 369 0 4.805e-15
c3646 397 290 1.58e-16
c3647 0 62 1.05e-15
c3648 113 135 1.88e-16
c3649 246 226 7.96e-16
c3650 298 1 1.327e-15
c3651 417 238 1.58e-16
c3652 28 27 7.32e-16
c3653 327 282 7.96e-16
c3654 3 44 1.58e-16
c3655 0 17 3.756e-15
c3656 109 1 3.077e-15
c3657 206 441 1.58e-16
c3658 98 260 1.58e-16
c3659 151 1 8.3e-16
c3660 269 440 5.03e-16
c3661 50 0 1.827e-15
c3662 320 113 1.58e-16
c3663 440 3 3.15e-16
c3664 0 482 8.06e-16
c3665 104 0 3.154e-15
c3666 386 373 3.15e-16
c3667 100 53 9.74e-16
c3668 98 85 4.6e-16
c3669 77 78 4.8e-16
c3670 167 144 3.15e-16
c3671 158 0 8.3e-16
c3672 132 216 7.96e-16
c3673 175 230 3.15e-16
c3674 420 311 3.15e-16
c3675 89 1 4.616e-15
c3676 57 167 2.62e-16
c3677 50 113 1.58e-16
c3678 287 330 3.15e-16
c3679 326 290 1.58e-16
c3680 133 1 5.001e-15
c3681 342 57 1.9e-16
c3682 282 300 3.15e-16
c3683 309 307 3.15e-16
c3684 506 83 6.06e-16
c3685 1 106 3.163e-15
c3686 397 304 3.15e-16
c3687 143 0 7.35e-15
c3688 98 100 9.21e-16
c3689 140 39 7.32e-16
c3690 1 393 8.06e-16
c3691 464 459 1.132e-15
c3692 225 320 1.58e-16
c3693 320 30 1.74e-16
c3694 348 0 1.862e-15
c3695 381 386 3.54e-16
c3696 397 395 5.11e-16
c3697 142 114 3.15e-16
c3698 177 171 7.96e-16
c3699 271 272 3.306e-15
c3700 219 324 1.58e-16
c3701 225 306 1.58e-16
c3702 109 1 6.478e-15
c3703 260 181 1.58e-16
c3704 378 377 4.6e-16
c3705 363 1 4.427e-15
c3706 137 227 1.58e-16
c3707 135 28 9.74e-16
c3708 441 110 1.58e-16
c3709 50 30 1.58e-16
c3710 418 348 1.58e-16
c3711 4 5 1.88e-15
c3712 320 28 1.58e-16
c3713 1 149 7.665e-15
c3714 299 15 1.58e-16
c3715 1 438 1.565e-15
c3716 310 231 6.06e-16
c3717 502 411 1.58e-16
c3718 0 498 3.189e-15
c3719 413 513 1.042e-15
c3720 306 1 8.3e-16
c3721 397 464 1.58e-16
c3722 437 407 3.15e-16
c3723 1 503 3.163e-15
c3724 143 155 3.15e-16
c3725 468 472 1.6e-16
c3726 104 102 1.58e-16
c3727 269 364 6.3e-16
c3728 432 288 3.15e-16
c3729 96 164 1.58e-16
c3730 109 234 1.58e-16
c3731 100 181 4.73e-16
c3732 0 348 2.493e-15
c3733 226 164 1.58e-16
c3734 143 0 1.892e-15
c3735 231 303 9.74e-16
c3736 359 1 1.565e-15
c3737 124 0 1.827e-15
c3738 219 0 8.3e-16
c3739 449 1 3.293e-15
c3740 175 320 4.27e-16
c3741 145 114 1.58e-16
c3742 162 353 3.15e-16
c3743 451 395 3.306e-15
c3744 256 230 3.15e-16
c3745 420 503 3.15e-16
c3746 437 70 1.58e-16
c3747 76 53 1.58e-16
c3748 311 304 1.58e-16
c3749 369 476 1.58e-16
c3750 124 121 5.11e-16
c3751 491 238 6.62e-16
c3752 502 516 5.38e-16
c3753 294 299 3.15e-16
c3754 81 114 1.58e-16
c3755 512 415 3.137e-15
c3756 116 115 7.32e-16
c3757 149 1 2.565e-15
c3758 57 0 8.3e-16
c3759 70 161 1.58e-16
c3760 395 396 1.6e-16
c3761 357 347 1.58e-16
c3762 334 0 8.06e-16
c3763 401 332 7.96e-16
c3764 397 409 4.73e-16
c3765 200 197 1.042e-15
c3766 290 0 1.892e-15
c3767 420 0 1.05e-15
c3768 319 223 3.15e-16
c3769 271 113 7.32e-16
c3770 7 1 4.109e-15
c3771 19 0 3.055e-15
c3772 384 0 1.327e-15
c3773 363 373 1.58e-16
c3774 137 133 1.03e-16
c3775 226 15 1.58e-16
c3776 181 361 6.36e-16
c3777 130 129 6.36e-16
c3778 174 0 8.06e-16
c3779 316 397 4.73e-16
c3780 158 161 1.58e-16
c3781 385 386 1.03e-16
c3782 1 456 8.06e-16
c3783 106 108 1.926e-15
c3784 78 1 1.2359e-14
c3785 210 294 4.39e-16
c3786 0 291 2.493e-15
c3787 1 295 4.761e-15
c3788 134 0 8.06e-16
c3789 234 149 1.58e-16
c3790 250 1 8.3e-16
c3791 437 332 1.58e-16
c3792 57 155 1.58e-16
c3793 83 353 2.46e-16
c3794 326 1 2.565e-15
c3795 505 490 1.58e-16
c3796 0 144 3.306e-15
c3797 316 250 1.58e-16
c3798 0 488 2.912e-15
c3799 322 271 7.96e-16
c3800 219 281 1.58e-16
c3801 285 267 1.58e-16
c3802 295 114 1.58e-16
c3803 1 429 5.319e-15
c3804 96 65 1.58e-16
c3805 57 0 8.3e-16
c3806 304 0 1.892e-15
c3807 290 0 8.3e-16
c3808 295 207 1.58e-16
c3809 416 417 1.132e-15
c3810 55 78 1.58e-16
c3811 354 352 3.306e-15
c3812 24 300 1.58e-16
c3813 256 320 1.58e-16
c3814 1 267 3.724e-15
c3815 441 362 1.58e-16
c3816 124 300 1.58e-16
c3817 366 274 3.54e-16
c3818 30 46 1.58e-16
c3819 27 25 3.31e-16
c3820 115 107 1.58e-16
c3821 1 241 3.163e-15
c3822 252 149 9.54e-16
c3823 0 445 5.051e-15
c3824 169 114 1.58e-16
c3825 19 0 1.612e-15
c3826 418 304 1.58e-16
c3827 391 298 1.926e-15
c3829 1 433 1.565e-15
c3830 48 46 1.58e-16
c3831 75 0 3.724e-15
c3832 218 135 6.62e-16
c3833 311 1 1.327e-15
c3834 366 192 1.58e-16
c3835 170 166 1.58e-16
c3836 502 500 1.58e-16
c3837 432 287 3.15e-16
c3838 96 387 1.58e-16
c3839 113 19 1.58e-16
c3840 56 0 2.893e-15
c3841 28 46 3.15e-16
c3842 1 208 1.565e-15
c3843 0 167 1.612e-15
c3844 111 1 8.3e-16
c3845 1 30 3.163e-15
c3846 144 148 7.96e-16
c3847 331 299 7.96e-16
c3848 1 476 4.591e-15
c3849 0 304 4.427e-15
c3850 144 30 1.58e-16
c3851 354 1 1.565e-15
c3852 339 417 5.74e-16
c3853 96 53 3.15e-16
c3854 518 0 1.327e-15
c3855 100 1 2.514e-15
c3856 98 522 7.96e-16
c3857 0 465 8.06e-16
c3858 48 1 2.565e-15
c3859 0 395 2.476e-15
c3860 1 447 8.29e-15
c3861 294 105 1.58e-16
c3862 0 352 4.462e-15
c3863 28 134 7.96e-16
c3864 188 196 6.62e-16
c3865 48 144 1.58e-16
c3866 28 1 4.427e-15
c3867 418 214 1.58e-16
c3869 413 502 5.11e-16
c3870 28 144 3.15e-16
c3871 282 299 3.15e-16
c3872 420 476 3.15e-16
c3873 19 30 3.15e-16
c3874 319 193 3.15e-16
c3875 250 315 1.58e-16
c3876 109 162 1.58e-16
c3877 0 370 3.154e-15
c3878 100 420 1.58e-16
c3879 98 96 9.38e-16
c3880 155 167 1.58e-16
c3881 1 57 3.289e-15
c3882 0 32 3.756e-15
c3883 407 247 7.75e-16
c3884 8 10 1.926e-15
c3885 320 25 1.58e-16
c3886 169 173 1.58e-16
c3887 19 48 1.58e-16
c3888 447 384 1.58e-16
c3889 0 196 2.893e-15
c3890 167 0 3.756e-15
c3891 485 488 6.62e-16
c3892 3 193 3.15e-16
c3893 1 235 3.163e-15
c3894 157 158 7.32e-16
c3895 78 89 3.54e-16
c3896 131 0 8.06e-16
c3897 50 203 7.79e-16
c3898 0 426 8.06e-16
c3899 0 188 2.912e-15
c3900 1 198 3.189e-15
c3901 113 167 1.58e-16
c3902 72 0 3.756e-15
c3903 71 1 3.724e-15
c3904 212 1 3.163e-15
c3905 250 184 3.54e-16
c3906 24 47 7.96e-16
c3907 316 0 1.892e-15
c3908 156 1 1.565e-15
c3909 132 226 1.58e-16
c3910 0 490 8.811e-15
c3911 510 512 6.36e-16
c3912 502 514 3.306e-15
c3913 1 161 8.354e-15
c3914 293 324 1.58e-16
c3915 418 1 8.3e-16
c3916 59 1 1.565e-15
c3917 40 0 3.306e-15
c3918 70 319 1.58e-16
c3919 169 184 1.58e-16
c3920 206 192 1.58e-16
c3921 316 418 1.58e-16
c3922 70 500 8.89e-16
c3923 314 307 1.926e-15
c3924 201 0 8.3e-16
c3925 1 435 4.591e-15
c3926 0 12 1.862e-15
c3927 318 0 4.575e-15
c3928 290 286 1.58e-16
c3929 493 487 1.58e-16
c3930 110 112 1.926e-15
c3931 217 214 3.15e-16
c3932 418 114 1.58e-16
c3933 0 468 4.303e-15
c3935 151 353 1.58e-16
c3936 83 109 1.58e-16
c3937 109 283 1.58e-16
c3938 441 192 1.58e-16
c3939 0 409 5.898e-15
c3940 437 505 3.15e-16
c3941 295 116 1.58e-16
c3942 440 0 8.3e-16
c3943 342 313 1.58e-16
c3944 347 343 2.02e-16
c3945 136 34 1.042e-15
c3946 358 1 8.3e-16
c3947 0 443 3.194e-15
c3948 35 39 1.59e-15
c3949 86 1 1.862e-15
c3950 318 418 3.15e-16
c3951 342 225 3.15e-16
c3952 437 392 1.66e-16
c3953 96 369 1.58e-16
c3954 99 53 7.96e-16
c3955 316 0 8.3e-16
c3956 520 1 1.565e-15
c3957 125 107 3.54e-16
c3958 323 0 8.06e-16
c3959 219 151 6.3e-16
c3960 357 468 1.58e-16
c3961 0 495 8.06e-16
c3962 129 114 3.15e-16
c3963 264 101 6.36e-16
c3964 227 27 1.58e-16
c3965 40 54 7.96e-16
c3966 330 295 3.15e-16
c3967 158 159 2.038e-15
c3968 201 0 8.3e-16
c3969 342 1 8.3e-16
c3970 295 223 1.58e-16
c3971 164 39 1.58e-16
c3972 151 227 3.15e-16
c3973 318 0 3.223e-15
c3974 155 0 1.892e-15
c3975 231 319 3.15e-16
c3976 326 330 1.58e-16
c3977 447 395 2.6e-16
c3978 518 519 2.69e-15
c3979 234 235 7.32e-16
c3980 0 440 8.3e-16
c3981 1 157 2.247e-15
c3982 0 173 3.689e-15
c3983 86 88 3.306e-15
c3984 324 288 1.58e-16
c3985 352 85 1.58e-16
c3986 90 94 5.11e-16
c3987 95 1 3.083e-15
c3988 274 276 1.926e-15
c3989 0 315 2.493e-15
c3990 1 300 4.761e-15
c3991 436 409 6.62e-16
c3992 392 474 6.36e-16
c3993 64 0 1.05e-15
c3994 1 9 4.761e-15
c3995 256 57 1.58e-16
c3996 1 415 5.562e-15
c3997 175 167 2.62e-16
c3998 464 476 1.58e-16
c3999 432 390 1.58e-16
c4000 490 83 4.48e-16
c4001 509 506 7.96e-16
c4002 469 470 1.6e-16
c4003 0 486 3.154e-15
c4004 113 0 8.3e-16
c4005 353 62 1.58e-16
c4006 300 114 1.58e-16
c4007 295 107 1.58e-16
c4008 0 45 8.06e-16
c4009 219 363 1.58e-16
c4010 122 121 6.36e-16
c4011 300 207 1.58e-16
c4012 357 344 4.73e-16
c4013 24 299 1.58e-16
c4014 247 1 2.565e-15
c4015 219 320 1.58e-16
c4016 371 330 1.275e-15
c4017 420 415 3.15e-16
c4018 502 397 4.73e-16
c4019 15 39 3.15e-16
c4020 261 0 2.683e-15
c4021 124 299 2.62e-16
c4022 260 1 8.3e-16
c4023 135 227 1.88e-16
c4024 155 0 2.6e-15
c4025 332 298 3.15e-16
c4026 493 397 3.15e-16
c4027 432 487 3.15e-16
c4028 441 294 1.58e-16
c4029 319 1 8.3e-16
c4030 11 4 7.96e-16
c4031 320 227 1.58e-16
c4032 163 114 3.15e-16
c4033 157 1 4.616e-15
c4034 83 0 1.327e-15
c4035 283 0 8.3e-16
c4037 225 0 1.892e-15
c4038 1 504 8.06e-16
c4039 397 481 3.15e-16
c4040 1 115 3.724e-15
c4041 114 85 1.58e-16
c4042 1 25 6.864e-15
c4043 269 275 3.15e-16
c4044 3 1 2.247e-15
c4045 100 1 3.7e-15
c4046 113 0 3.194e-15
c4047 0 48 2.887e-15
c4048 162 241 1.263e-15
c4049 356 0 2.893e-15
c4050 437 0 8.3e-16
c4051 96 1 8.3e-16
c4052 38 36 1.926e-15
c4053 0 364 1.612e-15
c4054 497 498 2.69e-15
c4055 1 286 4.616e-15
c4056 326 481 4.48e-16
c4057 294 110 1.58e-16
c4058 517 516 6.62e-16
c4059 109 168 1.926e-15
c4060 256 167 3.15e-16
c4061 319 1 8.3e-16
c4062 151 109 1.58e-16
c4063 330 0 1.327e-15
c4064 397 407 3.15e-16
c4065 256 342 1.58e-16
c4066 357 437 1.58e-16
c4067 19 203 1.275e-15
c4068 342 381 3.15e-16
c4069 0 148 8.06e-16
c4070 0 223 1.444e-15
c4071 417 164 1.58e-16
c4072 432 459 1.58e-16
c4073 0 111 3.756e-15
c4074 175 0 4.006e-15
c4075 493 311 1.328e-15
c4076 115 1 1.327e-15
c4077 288 281 1.421e-15
c4078 488 306 1.58e-16
c4079 0 474 2.893e-15
c4080 287 324 1.58e-16
c4081 39 53 1.59e-15
c4082 3 1 3.289e-15
c4083 418 223 1.58e-16
c4084 1 361 3.083e-15
c4085 1 238 6.214e-15
c4086 90 87 3.15e-16
c4087 48 0 8.3e-16
c4088 159 1 4.761e-15
c4089 260 173 1.58e-16
c4090 70 397 4.73e-16
c4091 0 102 2.661e-15
c4092 215 0 8.06e-16
c4093 441 4 1.58e-16
c4094 440 5 1.58e-16
c4095 1 279 6.355e-15
c4096 28 0 5.551e-15
c4097 0 411 2.476e-15
c4098 113 48 3.15e-16
c4099 14 1 5.079e-15
c4100 0 330 1.444e-15
c4101 96 290 4.11e-16
c4102 432 397 1.58e-16
c4103 505 500 3.15e-16
c4104 1 489 1.565e-15
c4105 70 250 1.58e-16
c4106 219 267 1.58e-16
c4107 420 238 3.15e-16
c4108 417 15 1.58e-16
c4109 0 287 1.862e-15
c4110 100 173 1.58e-16
c4111 121 107 3.15e-16
c4112 260 184 3.54e-16
c4113 262 184 4.8e-16
c4114 56 58 6.36e-16
c4115 175 0 1.327e-15
c4116 452 373 6.36e-16
c4117 109 320 1.58e-16
c4118 357 411 3.15e-16
c4119 437 83 1.58e-16
c4120 111 30 3.15e-16
c4121 300 116 1.58e-16
c4122 86 0 1.892e-15
c4123 151 149 3.15e-16
VCin 193 0 pwl (0 0 8e-08 0 8.2e-08 3 1.6e-07 3 
+ 1.62e-07 0 )
VAin20 353 0 pwl (0 0 4e-08 0 4.2e-08 3 8e-08 3 
+ 8.2e-08 0 1.2e-07 0 1.22e-07 3 1.6e-07 3 
+ 1.62e-07 0 )
VAin19 320 0 pwl (0 0 1.2e-07 0 1.22e-07 3 1.6e-07 3 
+ 1.62e-07 0 )
VAin18 418 0 pwl (0 0 4e-08 0 4.2e-08 3 8e-08 3 
+ 8.2e-08 0 1.2e-07 0 1.22e-07 3 1.6e-07 3 
+ 1.62e-07 0 )
VAin17 72 0 pwl (0 0 1.2e-07 0 1.22e-07 3 1.6e-07 3 
+ 1.62e-07 0 )
VAin16 227 0 pwl (0 0 1.2e-07 0 1.22e-07 3 1.6e-07 3 
+ 1.62e-07 0 )
VAin15 145 0 pwl (0 0 4e-08 0 4.2e-08 3 8e-08 3 
+ 8.2e-08 0 1.2e-07 0 1.22e-07 3 1.6e-07 3 
+ 1.62e-07 0 )
VAin14 159 0 pwl (0 0 1.2e-07 0 1.22e-07 3 1.6e-07 3 
+ 1.62e-07 0 )
VAin13 164 0 pwl (0 0 4e-08 0 4.2e-08 3 8e-08 3 
+ 8.2e-08 0 1.2e-07 0 1.22e-07 3 1.6e-07 3 
+ 1.62e-07 0 )
VAin12 17 0 pwl (0 0 4e-08 0 4.2e-08 3 8e-08 3 
+ 8.2e-08 0 1.2e-07 0 1.22e-07 3 1.6e-07 3 
+ 1.62e-07 0 )
VAin11 41 0 pwl (0 0 1.2e-07 0 1.22e-07 3 1.6e-07 3 
+ 1.62e-07 0 )
VAin10 37 0 pwl (0 0 4e-08 0 4.2e-08 3 8e-08 3 
+ 8.2e-08 0 1.2e-07 0 1.22e-07 3 1.6e-07 3 
+ 1.62e-07 0 )
VAin9 111 0 pwl (0 0 1.2e-07 0 1.22e-07 3 1.6e-07 3 
+ 1.62e-07 0 )
VAin8 441 0 pwl (0 0 1.2e-07 0 1.22e-07 3 1.6e-07 3 
+ 1.62e-07 0 )
VAin7 295 0 pwl (0 0 4e-08 0 4.2e-08 3 8e-08 3 
+ 8.2e-08 0 1.2e-07 0 1.22e-07 3 1.6e-07 3 
+ 1.62e-07 0 )
VAin6 283 0 pwl (0 0 1.2e-07 0 1.22e-07 3 1.6e-07 3 
+ 1.62e-07 0 )
VAin5 300 0 pwl (0 0 4e-08 0 4.2e-08 3 8e-08 3 
+ 8.2e-08 0 1.2e-07 0 1.22e-07 3 1.6e-07 3 
+ 1.62e-07 0 )
VAin4 5 0 pwl (0 0 4e-08 0 4.2e-08 3 8e-08 3 
+ 8.2e-08 0 1.2e-07 0 1.22e-07 3 1.6e-07 3 
+ 1.62e-07 0 )
VAin3 9 0 pwl (0 0 1.2e-07 0 1.22e-07 3 1.6e-07 3 
+ 1.62e-07 0 )
VAin2 32 0 pwl (0 0 4e-08 0 4.2e-08 3 8e-08 3 
+ 8.2e-08 0 1.2e-07 0 1.22e-07 3 1.6e-07 3 
+ 1.62e-07 0 )
VAin1 21 0 pwl (0 0 1.2e-07 0 1.22e-07 3 1.6e-07 3 
+ 1.62e-07 0 )
VBin20 352 0 pwl (0 0 8e-08 0 8.2e-08 3 1.2e-07 3 
+ 1.22e-07 0 1.6e-07 0 )
VBin19 319 0 pwl (0 0 4e-08 0 4.2e-08 3 1.2e-07 3 
+ 1.22e-07 0 1.6e-07 0 )
VBin18 417 0 pwl (0 0 8e-08 0 8.2e-08 3 1.2e-07 3 
+ 1.22e-07 0 1.6e-07 0 )
VBin17 71 0 pwl (0 0 4e-08 0 4.2e-08 3 1.2e-07 3 
+ 1.22e-07 0 1.6e-07 0 )
VBin16 226 0 pwl (0 0 4e-08 0 4.2e-08 3 1.2e-07 3 
+ 1.22e-07 0 1.6e-07 0 )
VBin15 144 0 pwl (0 0 8e-08 0 8.2e-08 3 1.2e-07 3 
+ 1.22e-07 0 1.6e-07 0 )
VBin14 158 0 pwl (0 0 4e-08 0 4.2e-08 3 1.2e-07 3 
+ 1.22e-07 0 1.6e-07 0 )
VBin13 163 0 pwl (0 0 8e-08 0 8.2e-08 3 1.2e-07 3 
+ 1.22e-07 0 1.6e-07 0 )
VBin12 16 0 pwl (0 0 8e-08 0 8.2e-08 3 1.2e-07 3 
+ 1.22e-07 0 1.6e-07 0 )
VBin11 40 0 pwl (0 0 4e-08 0 4.2e-08 3 1.2e-07 3 
+ 1.22e-07 0 1.6e-07 0 )
VBin10 36 0 pwl (0 0 8e-08 0 8.2e-08 3 1.2e-07 3 
+ 1.22e-07 0 1.6e-07 0 )
VBin9 110 0 pwl (0 0 4e-08 0 4.2e-08 3 1.2e-07 3 
+ 1.22e-07 0 1.6e-07 0 )
VBin8 440 0 pwl (0 0 4e-08 0 4.2e-08 3 1.2e-07 3 
+ 1.22e-07 0 1.6e-07 0 )
VBin7 294 0 pwl (0 0 8e-08 0 8.2e-08 3 1.2e-07 3 
+ 1.22e-07 0 1.6e-07 0 )
VBin6 282 0 pwl (0 0 4e-08 0 4.2e-08 3 1.2e-07 3 
+ 1.22e-07 0 1.6e-07 0 )
VBin5 299 0 pwl (0 0 8e-08 0 8.2e-08 3 1.2e-07 3 
+ 1.22e-07 0 1.6e-07 0 )
VBin4 4 0 pwl (0 0 8e-08 0 8.2e-08 3 1.2e-07 3 
+ 1.22e-07 0 1.6e-07 0 )
VBin3 8 0 pwl (0 0 4e-08 0 4.2e-08 3 1.2e-07 3 
+ 1.22e-07 0 1.6e-07 0 )
VBin2 31 0 pwl (0 0 8e-08 0 8.2e-08 3 1.2e-07 3 
+ 1.22e-07 0 1.6e-07 0 )
VBin1 20 0 pwl (0 0 4e-08 0 4.2e-08 3 1.6e-07 3 
+ 1.62e-07 0 )
VVdd 1 0 3 
.temp 75 
.print TRAN v(342) v(437) v(518) v(497) v(432) v(420) 
+v(256) v(492) v(151) v(96) v(357) v(269) 
+v(449) v(467) v(458) v(475) v(201) v(285) 
+v(219) v(206) 
.options limpts=50000 itl5=50000
.TRAN 5e-10 1.6e-07
.end
